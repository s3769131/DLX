library ieee;
use ieee.std_logic_1164.all;
use work.CU_pkg.all;

entity cu_core is
  generic(
    CU_IR_NBIT : positive := 32);
  port(
    CU_instruction_register : in  std_logic_vector(CU_IR_NBIT - 1 downto 0);
    CU_decode_signed_ext    : out std_logic_vector(1 downto 0);
    CU_decode_dest_sel      : out std_logic_vector(1 downto 0);
    CU_decode_read1_en      : out std_logic;
    CU_decode_read2_en      : out std_logic;
    CU_execute_branch_type  : out std_logic;
    CU_execute_alu_op       : out std_logic_vector(5 downto 0);
    CU_execute_top_mux      : out std_logic;
    CU_execute_bottom_mux   : out std_logic;
    CU_execute_is_branch    : out std_logic;
    CU_memory_r_not_w       : out std_logic;
    CU_memory_signed_load   : out std_logic;
    CU_memory_load_type     : out std_logic_vector(1 downto 0);
    CU_writeback_write_en   : out std_logic;
    CU_writeback_mux        : out std_logic_vector(1 downto 0));
end entity;

architecture bhv of cu_core is
  signal s_cu_opcode : std_logic_vector(8 - 1 downto 0);
  signal s_cu_func   : std_logic_vector(8 - 1 downto 0);

begin
  s_cu_opcode(7 downto 6) <= (others => '0');
  s_cu_opcode(5 downto 0) <= CU_instruction_register(CU_IR_NBIT - 1 downto CU_IR_NBIT - CU_OPCODE_NBIT);
  
  s_cu_func(7 downto 6) <= (others => '0');
  s_cu_func(5 downto 0) <= CU_instruction_register(CU_FUNC_NBIT - 1 downto 0);

  MAIN : process(s_cu_opcode, s_cu_func)
  begin
    case (s_cu_opcode) is
      when CU_ALU_OPCODE =>
        case (s_cu_func) is
          when dlx_sll =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "001100"; --  sll
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_srl =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "000100"; --  srl
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_sra =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "000000"; --  sra
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_add =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "010000"; --  add
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_addu =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "010000"; --  add
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_sub =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "011000"; --  sub
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_subu =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "011000"; --  sub
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_and =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "111000"; --  and
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_or =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "111110"; --  or
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_xor =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "110110"; --  xor
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_seq =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "100100"; --  set equal
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_sne =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "100110"; --  set not equal
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_slt =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "100011"; --  set less than signed
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_sgt =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "101011"; --  set greater than signed
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_sle =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "100001"; --  set less equal signed
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_sge =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "101001"; --  set greater equal signed
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_sltu =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "100010"; --  set less than unsigned
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_sgtu =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "101010"; --  set greater than unsigned
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_sleu =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "100000"; --  set less equal unsigned
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when dlx_sgeu =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "10"; --  use rd as destination
            CU_decode_read1_en     <= '1'; --  read
            CU_decode_read2_en     <= '1'; --  read
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "101000"; --  set greater equal unsigned
            CU_execute_top_mux     <= '1'; --  take rs
            CU_execute_bottom_mux  <= '1'; --  take rt
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '1'; --  write to rf
            CU_writeback_mux       <= "01"; --  write data from ALU
          when others =>
            CU_decode_signed_ext   <= "00"; --  don't care
            CU_decode_dest_sel     <= "00"; --  write to 0
            CU_decode_read1_en     <= '0'; --  don't care
            CU_decode_read2_en     <= '0'; --  don't care
            CU_execute_branch_type <= '0'; --  don't care
            CU_execute_alu_op      <= "000000"; --  sll
            CU_execute_top_mux     <= '1'; --  don't care
            CU_execute_bottom_mux  <= '1'; --  don't care
            CU_execute_is_branch   <= '0'; --  is not branch
            CU_memory_r_not_w      <= '1'; --  don't write anything
            CU_memory_signed_load  <= '0'; --  don't care
            CU_memory_load_type    <= "00"; --  don't care
            CU_writeback_write_en  <= '0'; --  don't write to rf
            CU_writeback_mux       <= "00"; --  don't care
        end case;
      when dlx_j =>
        CU_decode_signed_ext   <= "01"; --  extend as 23 bits unsigned immediate
        CU_decode_dest_sel     <= "00"; --  don't care
        CU_decode_read1_en     <= '0';  --  don't read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '1';  --  j is always taken
        CU_execute_alu_op      <= "010000"; --  add immediate target to 0
        CU_execute_top_mux     <= '1';  --  read all zero from RF_in1
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '1';  --  is branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '0';  --  don't write anything
        CU_writeback_mux       <= "00"; --  don't care
      when dlx_jal =>
        CU_decode_signed_ext   <= "01"; --  extend as 23 bits unsigned immedaite
        CU_decode_dest_sel     <= "11"; --  force register 31 as destination
        CU_decode_read1_en     <= '0';  --  don't read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '1';  --  jal is always taken
        CU_execute_alu_op      <= "010000"; --  add immediate target to 0
        CU_execute_top_mux     <= '1';  --  read all zero from RF_in1
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '1';  --  is branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write npc to register 31
        CU_writeback_mux       <= "10"; --  write NPC
      when dlx_beqz =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immedaite
        CU_decode_dest_sel     <= "00"; --  don't care
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '1';  --  branch equal zero
        CU_execute_alu_op      <= "010000"; --  add
        CU_execute_top_mux     <= '0';  --  take NPC
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '1';  --  is branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '0';  --  don't write anything
        CU_writeback_mux       <= "00"; --  don't write anything
      when dlx_bnez =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immedaite
        CU_decode_dest_sel     <= "00"; --  don't care
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  branch not equal zero
        CU_execute_alu_op      <= "010000"; --  add
        CU_execute_top_mux     <= '0';  --  take NPC
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '1';  --  is branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '0';  --  don't write anything
        CU_writeback_mux       <= "00"; --  don't write anything
      when dlx_addi =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immedaite
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '1';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "010000"; --  add
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_addui =>
        CU_decode_signed_ext   <= "00"; --  extend as 16 bits unsigned immedaite
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '1';  --  read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "010000"; --  add
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_subi =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immedaite
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '1';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "011000"; --  sub
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_subui =>
        CU_decode_signed_ext   <= "00"; --  extend as 16 bits unsigned immedaite
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '1';  --  read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "011000"; --  sub
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_andi =>
        CU_decode_signed_ext   <= "00"; --  extend as 16 bits unsigned immedaite
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '1';  --  read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "111000"; --  and
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_ori =>
        CU_decode_signed_ext   <= "00"; --  extend as 16 bits unsigned immedaite
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '1';  --  read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "111110"; --  or
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_xori =>
        CU_decode_signed_ext   <= "00"; --  extend as 16 bits unsigned immedaite
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '1';  --  read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "110110"; --  xor
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      --when lhi    =>  --  still to do
      when dlx_jr =>
        CU_decode_signed_ext   <= "00"; --  don't care
        CU_decode_dest_sel     <= "00"; --  don't care
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '1';  --  absolute branch
        CU_execute_alu_op      <= "010000"; --  add
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  don't care
        CU_execute_is_branch   <= '1';  --  is branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '0';  --  don't write to rf
        CU_writeback_mux       <= "00"; --  don't care
      when dlx_jalr =>
        CU_decode_signed_ext   <= "00"; --  don't care
        CU_decode_dest_sel     <= "11"; --  force register 31 as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '1';  --  jalr is always taken
        CU_execute_alu_op      <= "010000"; --  add immediate target to 0
        CU_execute_top_mux     <= '1';  --  read rs
        CU_execute_bottom_mux  <= '1';  --  read all zero from RF_in2
        CU_execute_is_branch   <= '1';  --  is branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write npc to register 31
        CU_writeback_mux       <= "10"; --  write NPC
      when dlx_slli =>
        CU_decode_signed_ext   <= "00"; --  extend as 16 bits unsigned immedaite
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "001100"; --  sll
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_nop =>
        CU_decode_signed_ext   <= "00"; --  don't care
        CU_decode_dest_sel     <= "00"; --  write to 0
        CU_decode_read1_en     <= '0';  --  don't care
        CU_decode_read2_en     <= '0';  --  don't care
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "000000"; --  sll
        CU_execute_top_mux     <= '1';  --  don't care
        CU_execute_bottom_mux  <= '1';  --  don't care
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '0';  --  don't write to rf
        CU_writeback_mux       <= "00"; --  don't care
     
      when dlx_seqi =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "100100"; --  slt
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
        
        
        when dlx_snei =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "100110"; --  slt
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      
      
      when dlx_srli =>
        CU_decode_signed_ext   <= "00"; --  extend as 16 bits unsigned immedaite
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "000100"; --  srl
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_srai =>
        CU_decode_signed_ext   <= "00"; --  extend as 16 bits unsigned immedaite
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "000000"; --  sra
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_slti =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "100011"; --  slt
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_sgti =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "101011"; --  sgt
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_slei =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "100001"; --  sle
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_sgei =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "101001"; --  sge
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_lb =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "010000"; --  add
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  load
        CU_memory_signed_load  <= '1';  --  signed load
        CU_memory_load_type    <= "10"; --  load byte
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "00"; --  write data from MEM
      when dlx_lh =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "010000"; --  add
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  load
        CU_memory_signed_load  <= '1';  --  signed load
        CU_memory_load_type    <= "01"; --  load halfword
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "00"; --  write data from MEM
      when dlx_lw =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "010000"; --  add
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  load
        CU_memory_signed_load  <= '1';  --  signed load
        CU_memory_load_type    <= "00"; --  load word
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "00"; --  write data from MEM
      when dlx_lbu =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "010000"; --  add
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  load
        CU_memory_signed_load  <= '0';  --  unsigned load
        CU_memory_load_type    <= "10"; --  load byte
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "00"; --  write data from MEM
      when dlx_lhu =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "010000"; --  add
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  load
        CU_memory_signed_load  <= '0';  --  unsigned load
        CU_memory_load_type    <= "01"; --  load halfword
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "00"; --  write data from MEM
      when dlx_sw =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "010000"; --  add
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '0';  --  store
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "01"; --  don't care
        CU_writeback_write_en  <= '0';  --  don't write to rf
        CU_writeback_mux       <= "00"; --  don't   --  ?
      when dlx_sltui =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "100010"; --  slt
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_sgtui =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "101010"; --  sgt
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_sleui =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "100000"; --  sle
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when dlx_sgeui =>
        CU_decode_signed_ext   <= "10"; --  extend as 16 bits signed immediate
        CU_decode_dest_sel     <= "01"; --  use rt as destination
        CU_decode_read1_en     <= '1';  --  read
        CU_decode_read2_en     <= '0';  --  don't read
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "101000"; --  sge
        CU_execute_top_mux     <= '1';  --  take rs
        CU_execute_bottom_mux  <= '0';  --  read extended immediate from imm_in
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '1';  --  write to rf
        CU_writeback_mux       <= "01"; --  write data from ALU
      when others =>
        CU_decode_signed_ext   <= "00"; --  don't care
        CU_decode_dest_sel     <= "00"; --  write to 0
        CU_decode_read1_en     <= '0';  --  don't care
        CU_decode_read2_en     <= '0';  --  don't care
        CU_execute_branch_type <= '0';  --  don't care
        CU_execute_alu_op      <= "000000"; --  sll
        CU_execute_top_mux     <= '1';  --  don't care
        CU_execute_bottom_mux  <= '1';  --  don't care
        CU_execute_is_branch   <= '0';  --  is not branch
        CU_memory_r_not_w      <= '1';  --  don't write anything
        CU_memory_signed_load  <= '0';  --  don't care
        CU_memory_load_type    <= "00"; --  don't care
        CU_writeback_write_en  <= '0';  --  don't write to rf
        CU_writeback_mux       <= "00"; --  don't care
    end case;
  end process;

end architecture bhv;

configuration CFG_CU_CORE_BHV of cu_core is
  for bhv
  end for;
end configuration CFG_CU_CORE_BHV;
