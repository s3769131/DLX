package CONSTANTS is
  constant Nbit : integer := 32;
  constant Mbit : integer := 32;
end CONSTANTS;
