library ieee;
use ieee.std_logic_1164;

entity BTB is
  port (
    PC : in  std_logic_vector(31 downto 0);
    TARGET_PC :
    BRANCH_PREDICTION :
    CALCULATED_PC :
    CALCULATED_CONDITION :
    CLR
    EN
    RST
    CLK 
  );
end entity BTB;

architecture STR of BTB is

end architecture STR;
