
module DLX ( DLX_CLK, DLX_RST, ROM_ADDRESS, ROM_EN, ROM_DATA_READY, 
        ROM_INTERFACE, DRAM_ADDRESS, DRAM_EN, DRAM_READNOTWRITE, 
        DRAM_DATA_READY, DRAM_INTERFACE );
  output [31:0] ROM_ADDRESS;
  input [31:0] ROM_INTERFACE;
  output [31:0] DRAM_ADDRESS;
  inout [31:0] DRAM_INTERFACE;
  input DLX_CLK, DLX_RST, ROM_DATA_READY, DRAM_DATA_READY;
  output ROM_EN, DRAM_EN, DRAM_READNOTWRITE;
  wire   s_ID_rf_write_en, s_EX_IS_BRANCH, s_EX_BRANCH_TYPE, s_EX_BOT_MUX,
         s_MEM_SIGNED_LOAD,
         \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_up_network_p[1] ,
         \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_g[2] ,
         \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/CLA_PG_NET/N1 ,
         \core_inst/IF_stage/PLUS4_ADDER/RES_GENERATOR/CSA_15/sum_rca_0[1] ,
         \core_inst/IF_stage/PLUS4_ADDER/RES_GENERATOR/CSA_15/RCA_1/cout_tmp[0] ,
         \core_inst/IFID_NPC/DFF_3/N3 , \core_inst/IFID_NPC/DFF_5/N3 ,
         \core_inst/IFID_NPC/DFF_12/N3 , \core_inst/IFID_NPC/DFF_16/N3 ,
         \core_inst/IFID_IR/DFF_0/N3 , \core_inst/IFID_IR/DFF_1/N3 ,
         \core_inst/IFID_IR/DFF_3/N3 , \core_inst/IFID_IR/DFF_4/N3 ,
         \core_inst/IFID_IR/DFF_5/N3 , \core_inst/IFID_IR/DFF_6/N3 ,
         \core_inst/IFID_IR/DFF_7/N3 , \core_inst/IFID_IR/DFF_8/N3 ,
         \core_inst/IFID_IR/DFF_9/N3 , \core_inst/IFID_IR/DFF_10/N3 ,
         \core_inst/IFID_IR/DFF_11/N3 , \core_inst/IFID_IR/DFF_12/N3 ,
         \core_inst/IFID_IR/DFF_13/N3 , \core_inst/IFID_IR/DFF_14/N3 ,
         \core_inst/IFID_IR/DFF_15/N3 , \core_inst/IFID_IR/DFF_16/N3 ,
         \core_inst/IFID_IR/DFF_17/N3 , \core_inst/IFID_IR/DFF_18/N3 ,
         \core_inst/IFID_IR/DFF_19/N3 , \core_inst/IFID_IR/DFF_20/N3 ,
         \core_inst/IFID_IR/DFF_21/N3 , \core_inst/IFID_IR/DFF_22/N3 ,
         \core_inst/IFID_IR/DFF_23/N3 , \core_inst/IFID_IR/DFF_24/N3 ,
         \core_inst/IFID_IR/DFF_25/N3 , \core_inst/IFID_IR/DFF_26/N3 ,
         \core_inst/IFID_IR/DFF_27/N3 , \core_inst/IFID_IR/DFF_28/N3 ,
         \core_inst/IFID_IR/DFF_29/N3 , \core_inst/IFID_IR/DFF_30/N3 ,
         \core_inst/IFID_IR/DFF_31/N3 , \core_inst/IDEX_IR/DFF_26/N3 ,
         \core_inst/IDEX_IR/DFF_27/N3 , \core_inst/IDEX_IR/DFF_29/N3 ,
         \core_inst/IDEX_IR/DFF_30/N3 , \core_inst/IDEX_IR/DFF_31/N3 ,
         \core_inst/IDEX_NPC/DFF_0/N3 , \core_inst/IDEX_NPC/DFF_1/N3 ,
         \core_inst/IDEX_NPC/DFF_2/N3 , \core_inst/IDEX_NPC/DFF_3/N3 ,
         \core_inst/IDEX_NPC/DFF_4/N3 , \core_inst/IDEX_NPC/DFF_5/N3 ,
         \core_inst/IDEX_NPC/DFF_6/N3 , \core_inst/IDEX_NPC/DFF_7/N3 ,
         \core_inst/IDEX_NPC/DFF_8/N3 , \core_inst/IDEX_NPC/DFF_9/N3 ,
         \core_inst/IDEX_NPC/DFF_10/N3 , \core_inst/IDEX_NPC/DFF_11/N3 ,
         \core_inst/IDEX_NPC/DFF_12/N3 , \core_inst/IDEX_NPC/DFF_13/N3 ,
         \core_inst/IDEX_NPC/DFF_14/N3 , \core_inst/IDEX_NPC/DFF_15/N3 ,
         \core_inst/IDEX_NPC/DFF_16/N3 , \core_inst/IDEX_NPC/DFF_17/N3 ,
         \core_inst/IDEX_NPC/DFF_18/N3 , \core_inst/IDEX_NPC/DFF_19/N3 ,
         \core_inst/IDEX_NPC/DFF_20/N3 , \core_inst/IDEX_NPC/DFF_21/N3 ,
         \core_inst/IDEX_NPC/DFF_22/N3 , \core_inst/IDEX_NPC/DFF_24/N3 ,
         \core_inst/IDEX_NPC/DFF_25/N3 , \core_inst/IDEX_NPC/DFF_26/N3 ,
         \core_inst/IDEX_NPC/DFF_27/N3 , \core_inst/IDEX_NPC/DFF_28/N3 ,
         \core_inst/IDEX_NPC/DFF_29/N3 , \core_inst/IDEX_NPC/DFF_30/N3 ,
         \core_inst/IDEX_NPC/DFF_31/N3 , \core_inst/IDEX_RF_IN1/DFF_1/N3 ,
         \core_inst/IDEX_RF_IN1/DFF_2/N3 , \core_inst/IDEX_RF_IN1/DFF_3/N3 ,
         \core_inst/IDEX_RF_IN1/DFF_4/N3 , \core_inst/IDEX_RF_IN1/DFF_5/N3 ,
         \core_inst/IDEX_RF_IN1/DFF_6/N3 , \core_inst/IDEX_RF_IN1/DFF_7/N3 ,
         \core_inst/IDEX_RF_IN1/DFF_8/N3 , \core_inst/IDEX_RF_IN1/DFF_11/N3 ,
         \core_inst/IDEX_RF_IN1/DFF_12/N3 , \core_inst/IDEX_RF_IN1/DFF_13/N3 ,
         \core_inst/IDEX_RF_IN1/DFF_14/N3 , \core_inst/IDEX_RF_IN1/DFF_15/N3 ,
         \core_inst/IDEX_RF_IN1/DFF_19/N3 , \core_inst/IDEX_RF_IN1/DFF_20/N3 ,
         \core_inst/IDEX_RF_IN1/DFF_23/N3 , \core_inst/IDEX_RF_IN1/DFF_24/N3 ,
         \core_inst/IDEX_IMM_IN/DFF_0/N3 , \core_inst/IDEX_IMM_IN/DFF_1/N3 ,
         \core_inst/IDEX_IMM_IN/DFF_2/N3 , \core_inst/IDEX_IMM_IN/DFF_3/N3 ,
         \core_inst/IDEX_IMM_IN/DFF_4/N3 , \core_inst/IDEX_IMM_IN/DFF_5/N3 ,
         \core_inst/IDEX_IMM_IN/DFF_6/N3 , \core_inst/IDEX_IMM_IN/DFF_7/N3 ,
         \core_inst/IDEX_IMM_IN/DFF_8/N3 , \core_inst/IDEX_IMM_IN/DFF_9/N3 ,
         \core_inst/IDEX_IMM_IN/DFF_10/N3 , \core_inst/IDEX_IMM_IN/DFF_16/N3 ,
         \core_inst/IDEX_IMM_IN/DFF_17/N3 , \core_inst/IDEX_IMM_IN/DFF_18/N3 ,
         \core_inst/IDEX_IMM_IN/DFF_19/N3 , \core_inst/IDEX_IMM_IN/DFF_20/N3 ,
         \core_inst/IDEX_IMM_IN/DFF_21/N3 , \core_inst/IDEX_IMM_IN/DFF_22/N3 ,
         \core_inst/IDEX_IMM_IN/DFF_23/N3 , \core_inst/IDEX_IMM_IN/DFF_24/N3 ,
         \core_inst/IDEX_RF_IN2/DFF_0/N3 , \core_inst/IDEX_RF_IN2/DFF_1/N3 ,
         \core_inst/IDEX_RF_IN2/DFF_2/N3 , \core_inst/IDEX_RF_IN2/DFF_3/N3 ,
         \core_inst/IDEX_RF_IN2/DFF_4/N3 , \core_inst/IDEX_RF_IN2/DFF_5/N3 ,
         \core_inst/IDEX_RF_IN2/DFF_6/N3 , \core_inst/IDEX_RF_IN2/DFF_7/N3 ,
         \core_inst/IDEX_RF_IN2/DFF_8/N3 , \core_inst/IDEX_RF_IN2/DFF_13/N3 ,
         \core_inst/IDEX_RF_IN2/DFF_16/N3 , \core_inst/IDEX_RF_IN2/DFF_17/N3 ,
         \core_inst/IDEX_RF_IN2/DFF_18/N3 , \core_inst/IDEX_RF_IN2/DFF_19/N3 ,
         \core_inst/IDEX_RF_IN2/DFF_20/N3 , \core_inst/IDEX_RF_IN2/DFF_21/N3 ,
         \core_inst/IDEX_RF_IN2/DFF_23/N3 , \core_inst/IDEX_RF_IN2/DFF_24/N3 ,
         \core_inst/IDEX_RF_IN2/DFF_25/N3 , \core_inst/IDEX_RF_IN2/DFF_26/N3 ,
         \core_inst/IDEX_RF_IN2/DFF_27/N3 , \core_inst/IDEX_RF_IN2/DFF_28/N3 ,
         \core_inst/IDEX_RF_IN2/DFF_29/N3 ,
         \core_inst/IDEX_RF_ADDR_DEST/DFF_0/N3 ,
         \core_inst/IDEX_RF_ADDR_DEST/DFF_1/N3 ,
         \core_inst/IDEX_RF_ADDR_DEST/DFF_2/N3 ,
         \core_inst/IDEX_RF_ADDR_DEST/DFF_3/N3 ,
         \core_inst/IDEX_RF_ADDR_DEST/DFF_4/N3 ,
         \core_inst/EXMEM_IR/DFF_11/N3 , \core_inst/EXMEM_IR/DFF_12/N3 ,
         \core_inst/EXMEM_IR/DFF_13/N3 , \core_inst/EXMEM_IR/DFF_14/N3 ,
         \core_inst/EXMEM_IR/DFF_15/N3 , \core_inst/EXMEM_IR/DFF_16/N3 ,
         \core_inst/EXMEM_IR/DFF_17/N3 , \core_inst/EXMEM_IR/DFF_18/N3 ,
         \core_inst/EXMEM_IR/DFF_19/N3 , \core_inst/EXMEM_IR/DFF_20/N3 ,
         \core_inst/EXMEM_IR/DFF_26/N3 , \core_inst/EXMEM_IR/DFF_27/N3 ,
         \core_inst/EXMEM_IR/DFF_29/N3 , \core_inst/EXMEM_IR/DFF_30/N3 ,
         \core_inst/EXMEM_NPC/DFF_0/N3 , \core_inst/EXMEM_NPC/DFF_1/N3 ,
         \core_inst/EXMEM_NPC/DFF_2/N3 , \core_inst/EXMEM_NPC/DFF_3/N3 ,
         \core_inst/EXMEM_NPC/DFF_4/N3 , \core_inst/EXMEM_NPC/DFF_5/N3 ,
         \core_inst/EXMEM_NPC/DFF_6/N3 , \core_inst/EXMEM_NPC/DFF_7/N3 ,
         \core_inst/EXMEM_NPC/DFF_8/N3 , \core_inst/EXMEM_NPC/DFF_9/N3 ,
         \core_inst/EXMEM_NPC/DFF_10/N3 , \core_inst/EXMEM_NPC/DFF_11/N3 ,
         \core_inst/EXMEM_NPC/DFF_12/N3 , \core_inst/EXMEM_NPC/DFF_13/N3 ,
         \core_inst/EXMEM_NPC/DFF_14/N3 , \core_inst/EXMEM_NPC/DFF_15/N3 ,
         \core_inst/EXMEM_NPC/DFF_16/N3 , \core_inst/EXMEM_NPC/DFF_17/N3 ,
         \core_inst/EXMEM_NPC/DFF_18/N3 , \core_inst/EXMEM_NPC/DFF_19/N3 ,
         \core_inst/EXMEM_NPC/DFF_20/N3 , \core_inst/EXMEM_NPC/DFF_21/N3 ,
         \core_inst/EXMEM_NPC/DFF_22/N3 , \core_inst/EXMEM_NPC/DFF_23/N3 ,
         \core_inst/EXMEM_NPC/DFF_24/N3 , \core_inst/EXMEM_NPC/DFF_25/N3 ,
         \core_inst/EXMEM_NPC/DFF_26/N3 , \core_inst/EXMEM_NPC/DFF_27/N3 ,
         \core_inst/EXMEM_NPC/DFF_28/N3 , \core_inst/EXMEM_NPC/DFF_29/N3 ,
         \core_inst/EXMEM_NPC/DFF_30/N3 , \core_inst/EXMEM_NPC/DFF_31/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_0/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_1/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_2/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_3/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_4/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_5/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_6/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_7/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_8/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_9/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_10/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_11/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_12/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_13/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_14/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_15/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_16/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_17/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_18/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_19/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_20/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_21/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_22/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_23/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_24/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_25/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_26/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_27/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_28/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_29/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_30/N3 ,
         \core_inst/EXMEM_ALU_OUT/DFF_31/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_0/N3 , \core_inst/EXMEM_DATAIN/DFF_1/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_2/N3 , \core_inst/EXMEM_DATAIN/DFF_3/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_4/N3 , \core_inst/EXMEM_DATAIN/DFF_5/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_6/N3 , \core_inst/EXMEM_DATAIN/DFF_7/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_8/N3 , \core_inst/EXMEM_DATAIN/DFF_10/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_11/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_12/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_13/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_14/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_15/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_16/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_17/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_18/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_19/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_20/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_21/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_22/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_23/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_24/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_25/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_26/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_27/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_28/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_29/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_30/N3 ,
         \core_inst/EXMEM_DATAIN/DFF_31/N3 ,
         \core_inst/EXMEM_RF_ADDR_DEST/DFF_0/N3 ,
         \core_inst/EXMEM_RF_ADDR_DEST/DFF_1/N3 ,
         \core_inst/EXMEM_RF_ADDR_DEST/DFF_2/N3 ,
         \core_inst/EXMEM_RF_ADDR_DEST/DFF_3/N3 ,
         \core_inst/EXMEM_RF_ADDR_DEST/DFF_4/N3 ,
         \core_inst/MEMWB_IR/DFF_11/N3 , \core_inst/MEMWB_IR/DFF_12/N3 ,
         \core_inst/MEMWB_IR/DFF_13/N3 , \core_inst/MEMWB_IR/DFF_14/N3 ,
         \core_inst/MEMWB_IR/DFF_15/N3 , \core_inst/MEMWB_IR/DFF_16/N3 ,
         \core_inst/MEMWB_IR/DFF_17/N3 , \core_inst/MEMWB_IR/DFF_19/N3 ,
         \core_inst/MEMWB_IR/DFF_20/N3 , \core_inst/MEMWB_IR/DFF_30/N3 ,
         \core_inst/MEMWB_NPC/DFF_0/N3 , \core_inst/MEMWB_NPC/DFF_1/N3 ,
         \core_inst/MEMWB_NPC/DFF_2/N3 , \core_inst/MEMWB_NPC/DFF_3/N3 ,
         \core_inst/MEMWB_NPC/DFF_4/N3 , \core_inst/MEMWB_NPC/DFF_5/N3 ,
         \core_inst/MEMWB_NPC/DFF_6/N3 , \core_inst/MEMWB_NPC/DFF_7/N3 ,
         \core_inst/MEMWB_NPC/DFF_8/N3 , \core_inst/MEMWB_NPC/DFF_9/N3 ,
         \core_inst/MEMWB_NPC/DFF_10/N3 , \core_inst/MEMWB_NPC/DFF_11/N3 ,
         \core_inst/MEMWB_NPC/DFF_12/N3 , \core_inst/MEMWB_NPC/DFF_13/N3 ,
         \core_inst/MEMWB_NPC/DFF_14/N3 , \core_inst/MEMWB_NPC/DFF_15/N3 ,
         \core_inst/MEMWB_NPC/DFF_16/N3 , \core_inst/MEMWB_NPC/DFF_17/N3 ,
         \core_inst/MEMWB_NPC/DFF_18/N3 , \core_inst/MEMWB_NPC/DFF_19/N3 ,
         \core_inst/MEMWB_NPC/DFF_20/N3 , \core_inst/MEMWB_NPC/DFF_21/N3 ,
         \core_inst/MEMWB_NPC/DFF_22/N3 , \core_inst/MEMWB_NPC/DFF_23/N3 ,
         \core_inst/MEMWB_NPC/DFF_24/N3 , \core_inst/MEMWB_NPC/DFF_25/N3 ,
         \core_inst/MEMWB_NPC/DFF_26/N3 , \core_inst/MEMWB_NPC/DFF_27/N3 ,
         \core_inst/MEMWB_NPC/DFF_28/N3 , \core_inst/MEMWB_NPC/DFF_29/N3 ,
         \core_inst/MEMWB_NPC/DFF_30/N3 , \core_inst/MEMWB_NPC/DFF_31/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_0/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_1/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_2/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_3/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_4/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_5/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_6/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_7/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_8/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_9/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_10/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_11/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_12/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_13/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_14/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_15/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_16/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_17/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_18/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_19/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_20/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_21/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_22/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_23/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_24/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_25/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_26/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_27/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_28/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_29/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_30/N3 ,
         \core_inst/MEMWB_DATAOUT/DFF_31/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_0/N3 , \core_inst/MEMWB_ALUOUT/DFF_1/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_2/N3 , \core_inst/MEMWB_ALUOUT/DFF_3/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_4/N3 , \core_inst/MEMWB_ALUOUT/DFF_5/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_6/N3 , \core_inst/MEMWB_ALUOUT/DFF_7/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_8/N3 , \core_inst/MEMWB_ALUOUT/DFF_9/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_10/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_11/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_12/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_13/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_14/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_15/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_16/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_17/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_18/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_19/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_20/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_21/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_22/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_23/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_24/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_25/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_26/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_27/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_28/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_29/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_30/N3 ,
         \core_inst/MEMWB_ALUOUT/DFF_31/N3 ,
         \core_inst/MEMWB_RF_ADDR_DEST/DFF_0/N3 ,
         \core_inst/MEMWB_RF_ADDR_DEST/DFF_1/N3 ,
         \core_inst/MEMWB_RF_ADDR_DEST/DFF_2/N3 ,
         \core_inst/MEMWB_RF_ADDR_DEST/DFF_3/N3 ,
         \core_inst/MEMWB_RF_ADDR_DEST/DFF_4/N3 , \cu_inst/EX/DFF_1/N3 ,
         \cu_inst/EX/DFF_3/N3 , \cu_inst/EX/DFF_4/N3 , \cu_inst/EX/DFF_5/N3 ,
         \cu_inst/EX/DFF_6/N3 , \cu_inst/EX/DFF_7/N3 , \cu_inst/EX/DFF_9/N3 ,
         \cu_inst/EX/DFF_10/N3 , \cu_inst/EX/DFF_11/N3 ,
         \cu_inst/EX/DFF_12/N3 , \cu_inst/EX/DFF_13/N3 ,
         \cu_inst/EX/DFF_14/N3 , \cu_inst/EX/DFF_15/N3 ,
         \cu_inst/EX/DFF_16/N3 , \cu_inst/EX/DFF_17/N3 ,
         \cu_inst/EX/DFF_18/N3 , \cu_inst/MEM/DFF_0/N3 ,
         \cu_inst/MEM/DFF_1/N3 , \cu_inst/MEM/DFF_2/N3 ,
         \cu_inst/MEM/DFF_3/N3 , \cu_inst/MEM/DFF_4/N3 ,
         \cu_inst/MEM/DFF_5/N3 , \cu_inst/MEM/DFF_6/N3 , \cu_inst/WB/DFF_0/N3 ,
         \cu_inst/WB/DFF_1/N3 , \cu_inst/WB/DFF_2/N3 , \cu_inst/WB/DFF_3/N3 ,
         \core_inst/IF_stage/PROGRAM_COUNTER/DFF_0/N3 ,
         \core_inst/IF_stage/PROGRAM_COUNTER/DFF_1/N3 ,
         \core_inst/IF_stage/PROGRAM_COUNTER/DFF_2/N3 ,
         \core_inst/IF_stage/PROGRAM_COUNTER/DFF_10/N3 ,
         \core_inst/IF_stage/PROGRAM_COUNTER/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_1/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_2/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_3/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_4/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_5/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_6/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_7/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_8/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_9/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_10/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_11/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_12/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_13/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_14/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_15/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_16/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_17/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_18/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_19/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_20/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_21/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_22/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_23/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_24/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_25/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_26/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_27/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_28/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_29/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_30/DFF_31/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_0/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_1/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_2/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_3/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_4/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_5/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_6/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_7/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_8/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_9/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_10/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_11/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_12/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_13/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_14/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_15/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_16/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_17/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_18/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_19/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_20/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_21/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_22/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_23/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_24/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_25/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_26/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_27/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_28/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_29/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_30/N3 ,
         \core_inst/ID/REGISTER_FILE/REG_31/DFF_31/N3 ,
         \cu_inst/FW_UNIT/ITD_EXMEM/N17 , \cu_inst/FW_UNIT/ITD_EXMEM/N14 ,
         \core_inst/N65 , n297, n298, n334, n335, n336, n337, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n356, n358, n359, n360, n361, n363, n367, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n394, n396, n397, n398, n399,
         n401, n410, n411, n412, n413, n414, n415, n416, n417, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n432, n434,
         n435, n436, n437, n439, n446, n447, n448, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n461, n462, n463, n464, n465, n468,
         n469, n470, n471, n472, n473, n474, n475, n478, n482, n484, n485,
         n486, n487, n488, n489, n490, n491, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n506, n508, n509, n510, n511,
         n513, n522, n524, n525, n526, n527, n528, n529, n530, n531, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n546,
         n548, n549, n550, n551, n553, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n585, n587, n588, n589, n590, n592, n600,
         n602, n603, n604, n605, n606, n607, n608, n609, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n624, n626, n627,
         n628, n629, n631, n640, n642, n643, n644, n645, n646, n647, n648,
         n649, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n664, n666, n667, n668, n669, n671, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n703, n705, n706, n707, n708,
         n710, n716, n717, n719, n720, n721, n722, n723, n724, n725, n726,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n741, n743, n744, n745, n746, n748, n753, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n779, n781, n782, n783, n784,
         n786, n790, n793, n794, n796, n797, n798, n799, n800, n801, n802,
         n803, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n818, n820, n821, n822, n823, n825, n829, n834, n836, n837,
         n838, n839, n840, n841, n842, n843, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n858, n860, n861, n862, n863,
         n865, n869, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n897, n899, n900, n901, n902, n904, n912, n914, n915, n916,
         n917, n918, n919, n920, n921, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n936, n938, n939, n940, n941, n943,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n976,
         n978, n979, n980, n981, n983, n991, n993, n994, n995, n996, n997,
         n998, n1064, n1182, n1187, n1222, n1301, n1378, n1442, n1456, n1481,
         n1498, n1501, n1537, n1539, n1600, n1628, n1637, n1641, n1643, n1649,
         n1651, n1655, n1659, n1660, n1665, n1666, n1668, n1677, n1678, n1684,
         n1690, n1692, n1694, n1696, n1698, n1700, n1702, n1704, n1706, n1708,
         n1710, n1712, n1714, n1716, n1718, n1720, n1722, n1724, n1726, n1728,
         n1730, n1732, n1734, n1736, n1738, n1740, n1742, n1744, n1746, n1748,
         n1750, n1752, n1755, n2009, n2010, n2012, n2013, n2015, n2016, n2018,
         n2019, n2025, n2026, n2028, n2029, n2031, n2032, n2034, n2035, n2045,
         n2046, n2048, n2049, n2051, n2052, n2054, n2055, n2061, n2062, n2064,
         n2065, n2067, n2068, n2070, n2071, n2081, n2082, n2084, n2085, n2087,
         n2088, n2090, n2091, n2097, n2098, n2100, n2101, n2103, n2104, n2106,
         n2107, n2117, n2118, n2120, n2121, n2123, n2124, n2126, n2127, n2133,
         n2134, n2136, n2137, n2139, n2140, n2142, n2143, n2153, n2154, n2156,
         n2157, n2159, n2160, n2162, n2163, n2169, n2170, n2172, n2173, n2175,
         n2176, n2178, n2179, n2189, n2190, n2192, n2193, n2195, n2196, n2198,
         n2199, n2205, n2206, n2208, n2209, n2211, n2212, n2214, n2215, n2297,
         n2298, n2300, n2301, n2303, n2304, n2306, n2307, n2313, n2314, n2316,
         n2317, n2319, n2320, n2322, n2323, n2693, n2694, n2696, n2697, n2699,
         n2700, n2702, n2703, n2709, n2710, n2712, n2713, n2715, n2716, n2718,
         n2719, n2873, n2874, n2876, n2877, n2879, n2880, n2882, n2883, n2889,
         n2890, n2892, n2893, n2895, n2896, n2898, n2899, n2909, n2910, n2912,
         n2913, n2915, n2916, n2918, n2919, n2925, n2926, n2928, n2929, n2931,
         n2932, n2934, n2935, n2948, n2951, n2952, n2954, n2961, n2962, n2964,
         n2965, n2968, n2981, n2982, n2984, n2985, n2987, n2988, n2990, n2991,
         n2997, n2998, n3000, n3001, n3003, n3004, n3006, n3007, n3017, n3018,
         n3020, n3021, n3023, n3024, n3026, n3027, n3033, n3034, n3036, n3037,
         n3039, n3040, n3042, n3043, n3053, n3054, n3056, n3057, n3059, n3060,
         n3062, n3063, n3069, n3070, n3072, n3073, n3075, n3076, n3078, n3079,
         n3089, n3090, n3097, n3098, n3102, n3103, n3107, n3108, n3117, n3118,
         n3124, n3125, n3130, n3131, n3134, n3135, n4325, n4331, n4337, n4343,
         n4344, n4346, n4347, n4352, n4355, n4356, n4358, n4361, n4364, n4367,
         n4368, n4373, n4379, n4382, n4385, n4388, n4391, n4394, n4397, n4400,
         n4401, n4404, n4406, n4409, n4410, n4412, n4415, n4416, n4418, n4421,
         n4422, net81266, net89402, net89524, n5171, n5174, n5181, n5186,
         n5187, n5307, n5576, n5577, n5582, n5585, n5587, n5589, n5595, n5596,
         n5598, n5601, n5602, n5607, n5609, n5610, n5611, n5613, n5618, n5664,
         n5707, n5729, n5761, n6156, n6180, n6330, n6402, n6460, n6461, n6462,
         n6475, n6511, n6512, n6514, n6516, n6546, n6555, n6562, n6695, n6740,
         n6746, net334510, net342852, net342954, net342960, net342961,
         net342963, net365821, net365826, net366126, net366191, net366211,
         net366410, net366411, net366451, net366478, net366479, net366531,
         net399701, n11725, n11743, n11847, n11848, n11928, n13165, n13343,
         n13778, n13805, n13824, n14058, n14073, n14127, n14128, n14130,
         n14190, n14191, n14195, n14210, n14382, n14389, n14393, n14399,
         n14400, n14401, n14402, n14429, n14464, n14758, n14764, n14769,
         n15062, n15079, n16384, n16388, n16391, n17654, n17656, n17657,
         n17659, n17663, n17664, n17665, n17667, n17670, n17674, n17675,
         n17677, n17678, n17679, n17680, n17681, n17682, n17683, n17684,
         n17685, n17686, n17687, n17688, n17689, n17690, n17691, n17692,
         n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700,
         n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708,
         n17709, n17710, n17711, n17712, n17713, n17715, n17716, n17717,
         n17718, n17719, n17720, n17722, n17723, n17724, n17725, n17726,
         n17727, n17728, n17729, n17730, n17731, n17732, n17733, n17734,
         n17735, n17736, n17737, n17738, n17739, n17740, n17741, n17742,
         n17743, n17744, n17745, n17746, n17747, n17748, n17749, n17750,
         n17751, n17752, n17753, n17754, n17755, n17756, n17757, n17758,
         n17759, n17760, n17761, n17762, n17763, n17764, n17765, n17766,
         n17767, n17768, n17769, n17770, n17771, n17772, n17773, n17774,
         n17775, n17776, n17777, n17778, n17779, n17780, n17781, n17782,
         n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790,
         n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798,
         n17799, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17900, n17903, n17904, n17905, n17906, n17908, n17909, n17910,
         n17911, n17912, n17915, n17918, n17919, n17920, n17921, n17923,
         n17924, n17925, n17926, n17927, n17928, n17931, n17934, n17935,
         n17936, n17937, n17939, n17940, n17941, n17942, n17943, n17944,
         n17947, n17950, n17951, n17952, n17953, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17973, n17974,
         n17975, n17976, n17979, n17982, n17983, n17984, n17985, n17987,
         n17988, n17989, n17990, n17991, n17992, n17995, n17998, n17999,
         n18000, n18001, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18031, n18032, n18033, n18034, n18035, n18036,
         n18038, n18039, n18040, n18041, n18042, n18046, n18047, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18058, n18059,
         n18062, n18063, n18064, n18065, n18066, n18129, n18131, n18132,
         n18133, n18135, n18136, n18138, n18139, n18140, n18143, n18145,
         n18146, n18150, n18151, n18152, n18153, n18154, n18156, n18158,
         n18159, n18161, n18162, n18164, n18166, n18169, n18170, n18171,
         n18172, n18175, n18179, n18181, n18182, n18187, n18188, n18190,
         n18193, n18196, n18198, n18200, n18201, n18203, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18304, n18305, n18306,
         n18307, n18310, n18311, n18312, n18313, n18314, n18315, n18316,
         n18318, n18321, n18322, n18323, n18324, n18325, n18326, n18328,
         n18329, n18330, n18331, n18332, n18334, n18335, n18336, n18337,
         n18338, n18339, n18343, n18346, n18347, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18367, n18369, n18372, n18373,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18390, n18392, n18393, n18394, n18395, n18396, n18398,
         n18399, n18400, n18401, n18410, n18411, n18412, n18413, n18424,
         n18425, n18426, n18427, n18428, n18429, n18431, n18432, n18433,
         n18474, n18475, n18476, n18477, n18488, n18489, n18490, n18491,
         n18492, n18493, n18495, n18496, n18497, n18529, n18567, n18568,
         n18569, n18570, n18571, n18572, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18584, n18585, n18586, n18596,
         n18597, n18598, n18599, n18609, n18610, n18611, n18612, n18613,
         n18614, n18616, n18617, n18618, n18679, n18680, n18681, n18682,
         n18683, n18684, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18696, n18697, n18698, n18760, n18761, n18762,
         n18763, n18764, n18765, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18777, n18778, n18779, n18787, n18788,
         n18789, n18790, n18791, n18792, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18804, n18805, n18806, n18980,
         n18981, n18982, n18983, n18984, n18985, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18997, n18998, n18999,
         n19034, n19035, n19036, n19037, n19038, n19039, n19041, n19042,
         n19043, n19044, n19047, n19048, n19049, n19050, n19054, n19075,
         n19082, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19100, n19101, n19104, n19105, n19106, n19107, n19110,
         n19117, n19118, n19119, n19120, n19121, n19122, n19124, n19125,
         n19126, n19127, n19130, n19131, n19132, n19133, n19137, n19145,
         n19146, n19147, n19148, n19149, n19150, n19152, n19153, n19154,
         n19155, n19158, n19159, n19160, n19161, n19165, n19173, n19174,
         n19175, n19176, n19177, n19178, n19180, n19181, n19182, n19183,
         n19186, n19187, n19188, n19189, n19193, n19201, n19202, n19203,
         n19204, n19205, n19206, n19208, n19209, n19210, n19211, n19214,
         n19215, n19216, n19217, n19221, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19248, n19249, n19250, n19251, n19252,
         n19253, n19254, n19255, n19256, n19257, n19261, n19262, n19264,
         n19265, n19266, n19267, n19268, n19269, n19275, n19282, n19288,
         n19289, n19291, n19292, n19294, n19308, n19314, n19315, n19318,
         n19319, n19320, n19323, n19324, n19326, n19327, n19328, n19332,
         n19333, n19334, n19335, n19336, n19337, n19338, n19344, n19345,
         n19348, n19350, n19351, n19365, n19366, n19367, n19370, n19372,
         n19373, n19378, n19383, n19384, n19385, n19388, n19389, n19390,
         n19393, n19395, n19396, n19400, n19401, n19402, n19403, n19404,
         n19405, n19406, n19407, n19408, n19409, n19410, n19411, n19412,
         n19413, n19414, n19415, n19416, n19417, n19418, n19427, n19428,
         n19429, n19430, n19433, n19434, n19435, n19436, n19437, n19438,
         n19439, n19440, n19441, n19449, n19450, n19451, n19452, n19455,
         n19456, n19457, n19458, n19459, n19460, n19461, n19462, n19463,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19520, n19521, n19522, n19523, n19524, n19525, n19526, n19527,
         n19528, n19529, n19530, n19531, n19532, n19533, n19534, n19535,
         n19536, n19537, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19565, n19566, n19567,
         n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575,
         n19576, n19577, n19578, n19579, n19580, n19581, n19587, n19588,
         n19589, n19590, n19591, n19592, n19593, n19594, n19595, n19596,
         n19597, n19598, n19599, n19600, n19601, n19602, n19603, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638,
         n19639, n19640, n19641, n19642, n19643, n19644, n19645, n19646,
         n19647, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19773, n19774, n19775,
         n19776, n19777, n19778, n19779, n19787, n19788, n19789, n19790,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19851, n19852, n19853, n19854, n19855,
         n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863,
         n19864, n19865, n19866, n19867, n19873, n19874, n19875, n19876,
         n19877, n19878, n19879, n19880, n19881, n19882, n19883, n19884,
         n19885, n19886, n19887, n19888, n19889, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19952, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19969, n19970,
         n19971, n20011, n20012, n20013, n20041, n20042, n20049, n20054,
         n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062,
         n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070,
         n20071, n20072, n20073, n20074, n20075, n20076, n20077, n20078,
         n20080, n20081, n20084, n20085, n20086, n20087, n20088, n20092,
         n20107, n20110, n20111, n20117, n20118, n20134, n20153, n20154,
         n20155, n20182, n20183, n20200, n20201, n20202, n20204, n20220,
         n20221, n20223, n20240, n20241, n20243, n20260, n20261, n20263,
         n20293, n20294, n20296, n20313, n20315, n20332, n20333, n20334,
         n20350, n20351, n20367, n20368, n20370, n20371, n20372, n20373,
         n20375, n20392, n20394, n20396, n20397, n20398, n20400, n20431,
         n20432, n20433, n20443, n20445, n20462, n20464, n20481, n20483,
         n20501, n20502, n20519, n20521, n20547, n20549, n20581, n20582,
         n20592, n20593, n20609, n20610, n20611, n20613, n20630, n20632,
         n20650, n20651, n20667, n20668, n20684, n20686, n20704, n20706,
         net518455, net518461, net521855, net522736, net708964, net709330,
         net710357, net710387, net712313, net712344, net712353, net712356,
         net712365, net712377, net712378, net712384, net712390, net712391,
         net712397, net712445, net712462, net712466, net712467, net712468,
         net712469, net712472, net712488, net712490, net712493, net712494,
         net712499, net712520, net712606, net712737, net712795, net712808,
         net712812, net712838, net712847, net712855, net712856, net712857,
         net712872, net712879, net712880, net712882, net712886, net712893,
         net712922, net712931, net712945, net712961, net712971, net712975,
         net712976, net713148, net713151, net713152, net713154, net713167,
         net713168, net713389, net713412, net713414, net713438, net713442,
         net713448, net713454, net713463, net713467, net713468, net713554,
         net713560, net713561, net713564, net713570, net713602, net713606,
         net713607, net713612, net713627, net713633, net713636, net713669,
         net713672, net713677, net713679, net713681, net713683, net713687,
         net713692, net713701, net713707, net713711, net713726, net713728,
         net713736, net713738, net713740, net713748, net713751, net713753,
         net713754, net713760, net713761, net713762, net713763, net713767,
         net713770, net713773, net713777, net713779, net713785, net713810,
         net713811, net713829, net713845, net713849, net713850, net713857,
         net713863, net713866, net713867, net713868, net713869, net713870,
         net713873, net713874, net713882, net713892, net713894, net713897,
         net713905, net713906, net713907, net713923, net713924, net713930,
         net713934, net713949, net713950, net713951, net713952, net713964,
         net713967, net713977, net713978, net713979, net713985, net713990,
         net714006, net714007, net714033, net714034, net714076, net714077,
         net714104, net714105, net714113, net714122, net714123, net714157,
         net714164, net714182, net714194, net714249, net714251, net714261,
         net714267, net714275, net714281, net714287, net714306, net714309,
         net714335, net714344, net714346, net714347, net714354, net714378,
         net714382, net714401, net714440, net714463, net714464, net714465,
         net714466, net714486, net714487, net714488, net714489, net714494,
         net714542, net714544, net714551, net714559, net714585, net714602,
         net714603, net714611, net714612, net714751, net714754, net714756,
         net714770, net714845, net714855, net714858, net714861, net714871,
         net714877, net714907, net714934, net714943, net714965, net714977,
         net715015, net715018, net715019, net715027, net715032, net715048,
         net715058, net715169, net715170, net715175, net715200, net715221,
         net715235, net715284, net715313, net715359, net715419, net715420,
         net715421, net715422, net715443, net715460, net715584, net715586,
         net715591, net715592, net715614, net715632, net715656, net715661,
         net715668, net715705, net715706, net715707, net715794, net715795,
         net715796, net715842, net715847, net715884, net715885, net715892,
         net716231, net716223, net716221, net716215, net716237, net716369,
         net716367, net716353, net716341, net716337, net716333, net716331,
         net716313, net716311, net716267, net716261, net716259, net716255,
         net716249, net716247, net716243, net716387, net716405, net716417,
         net716423, net716461, net716477, net716491, net717048, net717050,
         net717049, net717052, net717053, net717056, net717055, net717060,
         net717074, net717087, net717091, net717106, net717105, net717104,
         net717103, net717153, net717157, net717454, net717463, net717511,
         net717510, net717547, net717570, net717720, net717719, net717718,
         net717789, net717830, net717843, net717876, net717875, net717926,
         net717952, net718006, net718033, net718070, net718069, net718074,
         net718078, net718077, net718081, net718082, net718087, net718086,
         net718092, net718098, net718103, net718111, net718134, net718133,
         net718139, net718138, net718152, net718154, net718337, net718341,
         net718340, net718349, net718351, net718355, net718361, net718367,
         net718372, net718380, net718391, net718400, net718405, net718432,
         net720121, net720303, n18972, n18971, n18970, n18964, n18860, n18859,
         n18858, n18855, n18854, n18853, n18852, n18851, n18850, n18849,
         n18848, n18846, n18845, n18844, n18843, n18842, n18841, n18644,
         n18643, n18642, n18639, n18638, n18637, n18636, n18635, n18634,
         n18633, n18632, n18630, n18629, n18628, n18627, n18626, n18625,
         n19929, n19928, n19927, n19925, n19924, n19923, n19922, n19921,
         n19920, n19919, n19918, n19917, n19916, n18725, n18724, n18723,
         n18720, n18719, n18718, n18717, n18716, n18715, n18714, n18713,
         n18711, n18710, n18709, n18708, n18707, n18706, net716385, n19394,
         n19391, n19387, n19382, n19381, n19380, n19379, n19377, n19376,
         n19375, n19374, n19364, n19363, n19362, n19361, n19360, n19359,
         n19358, n19357, n19493, n19490, n19489, n19485, n19484, n19483,
         n19482, n19479, n19478, n19476, n19475, n19474, n19473, n19472,
         n19470, n19469, net724632, net724631, net724630, net715700, net725586,
         net725577, net725613, net714175, net714174, net714173, net714172,
         net714394, net726961, net726959, net715551, net728159, net728158,
         net728314, net728481, net728823, net729186, net713813, net713833,
         net730300, net714241, net714240, net714239, net713851, net731329,
         net731327, net731344, net731713, net714689, net715615, net732762,
         net732754, net732750, net733097, net714657, net717059, net713864,
         net733611, net714873, net714476, net734022, net734282, net734346,
         net734385, net734607, net735179, net717075, net712470, net717462,
         net736739, net737672, net737706, net737713, net713733, net737907,
         net738443, net738474, net738517, net738840, net739078, net739130,
         net715236, net717615, net740075, net714860, net740493, net740492,
         net740526, net715769, net740632, net740634, net740645, net740649,
         net740655, net740661, net740674, net740706, net740710, net740717,
         net740721, net740739, net740741, net740801, net740803, net740818,
         net740820, net740834, net740836, net740858, net740860, net740886,
         net740888, net740918, net740920, net740936, net740938, net740970,
         net740972, net740989, net740991, net741006, net741008, net741037,
         net741039, net741054, net741056, net741078, net741080, net741108,
         net741110, net741130, net741132, net741147, net741149, net741170,
         net741172, net741196, net741198, net741214, net741216, net741237,
         net741262, net741279, net741280, net741282, net741293, net741301,
         net741305, net741306, net741307, net741329, net741339, net741345,
         net741353, net741384, net741385, net741388, net741389, net741397,
         net741400, net741440, net741442, net741456, net741458, net741464,
         net741518, net741520, net741525, net741527, net741531, net741532,
         net741539, net741541, net741544, net741547, net741549, net741565,
         net741572, net741576, net741580, net741582, net741603, net741608,
         net741609, net741620, net741686, net741696, net741726, net741959,
         net741958, net741987, net741999, net742011, net742017, net742037,
         net742042, net742047, net742046, net742061, net742087, net742092,
         net742100, net742146, net742157, net742182, net742198, net742209,
         net742224, net742243, net742242, net742241, net742248, net742259,
         net742265, net742271, net742275, net742286, net742284, net742296,
         net742304, net742309, net742315, net742326, net742325, net742324,
         net742331, net742339, net742368, net742413, net742412, net742423,
         net742473, net742483, net742508, net742507, net742506, net742593,
         net742649, net713208, net740076, n18752, n18751, n18750, n18747,
         n18746, n18745, n18744, n18743, n18742, n18741, n18740, n18738,
         n18737, n18736, n18735, n18734, n18733, n18945, n18944, n18943,
         n18940, n18939, n18938, n18937, n18936, n18935, n18934, n18933,
         n18931, n18930, n18929, n18928, n18927, n18926, net716257, net746701,
         net746688, net746687, net746753, net715020, net747343, net747437,
         net748275, net748274, net748269, net747347, net717543, net737101,
         net732533, net715647, net749230, net749260, net749274, net749273,
         net749289, net749292, net749295, net749308, net749307, net749306,
         net749312, net749317, net749334, net749338, net749343, net749363,
         net749369, net749372, net749375, net749387, net749408, net749410,
         net749427, net749428, net749439, net749434, net749443, net749442,
         net749454, net749465, net749476, net749489, net749495, net749507,
         net749525, net749529, net749533, net749534, net749542, net749551,
         net749566, net749612, net749636, net749664, net749679, net749685,
         net749698, net749697, net749707, net749710, net749709, net749725,
         net749732, net749798, net749806, net749812, net749817, net749823,
         net749822, net749820, net749830, net749832, net749841, net749843,
         net749894, net749898, net749905, net749910, net749922, net749926,
         net749930, net749936, net749945, net749951, net749967, net749972,
         net749977, net749987, net749993, net750019, net750025, net750024,
         net750032, net750053, net750057, net750086, net750090, net750093,
         net750135, net750158, net750176, net750182, net750203, net750228,
         net750238, net750255, net750264, net750274, net750277, net750278,
         net750287, net750290, net742612, net749902, net749500, net749839,
         net736366, net736356, net715528, net746315, net714508, net714507,
         net714506, net717845, net718083, net754762, net754997, net755033,
         net755048, net755056, net755060, net755061, net755075, net755086,
         net755090, net755097, net755134, net755137, net755139, net755207,
         net755210, net755214, net755216, net755238, net755241, net755240,
         net755255, net755258, net755260, net755610, net755637, net755683,
         net755699, net755708, net755714, net755733, net755740, net755757,
         net755745, net740679, net731199, net725127, net725126, net720370,
         net720369, net720368, net714575, net714553, net714552, net758037,
         net750122, net715666, net758544, net728824, net758644, net753553,
         net717461, net742223, net715445, net742012, net715672, net760144,
         net760161, net760170, n19910, n19908, n19907, n19906, n19905, n19904,
         n19903, n19902, n19901, n19900, n19899, n19898, n19897, n19896,
         n19895, net762579, net762597, net762604, net762625, net762654,
         net762661, net762660, net762674, net762729, net762754, net762753,
         net762759, net762762, n19994, n19992, n19991, n19990, n19989, n19988,
         n19987, n19986, n19985, n19984, n19983, n19982, n19981, n19980,
         n19979, n20036, n20034, n20033, n20032, n20031, n20030, n20029,
         n20028, n20027, n20026, n20025, n20024, n20023, n20022, n20021,
         net715662, net716263, net714975, net750085, net765319, net765341,
         net765340, net765429, net765546, net765629, net765727, net765730,
         net765744, net766652, net742648, net714610, net767167, net767168,
         net767169, net767171, net767172, net767173, net767203, net767205,
         net767206, net767207, net767208, net767209, net767210, net767211,
         net767214, net767221, net767232, net767234, net767235, net767237,
         net767238, net767239, net767257, net767320, net767330, net767335,
         net767341, net767340, net767352, net767357, net749400, net713806,
         net713805, net713804, net713803, net714947, net714724, net712473,
         net765361, net769908, net714749, net713710, net715176, net762680,
         net717760, net717742, \core_inst/EXMEM_IR/DFF_31/data_reg/n15 ,
         net715772, net715747, net750145, net713480, net773963, net773962,
         net773961, net738839, net724913, net724910, net765400, net714948,
         net715669, net762761, net762673, net714547, net714545, net714539,
         net714533, net714532, net714531, net714530, net714529, net758890,
         net749558, net714950, net715773, net755735, net742068, net714746,
         net729284, net714096, net733283, net733282, net715576, net715575,
         net714709, net714599, net737937, net762717, net766153, net715598,
         net745868, net745867, net742492, net755783, net714337, net713469,
         net745684, net745681, net745679, net745672, net714016, net749720,
         net718024, net748264, net750079, net742282, net715524, net740639,
         net717780, net717779, net717778, net715333, net729185, net729177,
         net715834, net737707, net714140, net715695, net729292, net729291,
         net750111, net715536, net715050, net715784, net715783, net755013,
         net769389, net768639, net714586, net713966, net755228, net750031,
         net736610, net736609, net763705, net714502, net714501, net712794,
         net712793, net715180, net755631, net715418, net720304, net720302,
         net729531, net729530, net725022, net713496, net713495, net715173,
         net765677, net713614, net715172, net715171, net714356, net714355,
         net714106, net778057, net778056, net778055, net755105, net715351,
         net712965, net713854, net755040, net778368, net714729, net724354,
         net724353, net724352, net733229, net733227, net778669, net714631,
         net742436, net715241, net714491, net714490, net713860, net713859,
         net713858, net755005, net734121, net713775, net714228, net714227,
         net714493, net714492, net712968, net712967, net712964, net713993,
         net713910, net713446, net741975, net755052, net749719, net749607,
         net738518, net742518, net717696, net712809, net713439, n20119, n18219,
         n18206, n18215, n18212, n18217, n18210, n18214, n18204, n18208,
         n18202, n18218, n18220, n18209, n18213, n18207, n18211, n18216,
         n18205, n20105, n20100, n20108, n20109, n20114, n20113, n20133,
         n20044, n20043, net713425, net713424, n20045, n18225, n18199, n18197,
         n18224, n18221, n18222, n18223, n19293, n19290, n18148, n18180,
         n18178, n18177, n18174, n18173, n18168, n18167, n18165, n18160,
         n18157, n18155, n18142, n18141, n18186, net780182, net780186,
         net780188, net780214, net780262, net780293, net780291, net780298,
         net780337, net780340, net780360, net780522, net780528, net780532,
         net780537, net780543, net780551, net780556, net780566, net780568,
         net780579, net780578, net780584, net780598, net780602, net714434,
         net714433, net714432, net714431, net714415, net714414, net714413,
         net714410, net714409, net781609, net727843, net727834, net727833,
         net727832, net727831, net727830, net782764, net731060, net716253,
         net717967, net783470, net783467, net783466, net714706, net715365,
         net780582, net742084, net715799, net715721, net715692, net716377,
         net716265, net742576, n15091, net716339, net731685, net715021,
         net784220, net714389, net714388, net714387, net714386, net714380,
         net714379, net784601, net718406, net713853, net714248, net717844,
         net749316, net732423, net741980, net713844, net742257, net785220,
         net785219, net785239, net785255, net785270, net785319, net740704,
         net714911, net714910, net714909, net714732, net714622, n13082,
         net749219, net717684, net786066, net742247, net715555, net765318,
         net731393, net715014, net749886, net765428, net786821, net786824,
         net786837, net786841, net786844, net786852, net786856, net786867,
         net787528, net787526, net787518, net787516, net787514, net787512,
         net780215, net749239, net746686, net734493, net717950, net713992,
         net713976, net713975, net713974, net713973, net713909, net712810,
         net712797, net712459, net712376, net767213, net750235, net748854,
         net735738, net735737, net735736, net735735, net734492, net725077,
         net720372, net718140, net717591, net715146, net714842, net714748,
         net714747, net714744, net714743, net714439, net714285, net714128,
         net714119, net714008, net714002, net713995, net794712, net795259,
         net795273, net795568, net795962, net796014, net796114, net796122,
         net796127, net796126, net796137, net796136, net796143, net796156,
         net796159, net796193, net796200, net796204, net796212, net796232,
         net796255, net796258, net796271, net795993, net780181, net713485,
         net713484, n20115, n18137, n18130, net749829, net720730, net720729,
         net720728, net720725, net720724, net715790, net715788, net804458,
         net804592, net804641, net804675, net804677, net796133, net785249,
         net780542, net780201, net780200, net755094, net738766, net738751,
         net736102, net726730, net726729, net713943, net713758, net713757,
         net713756, net713755, net713494, net713493, net713492, net713074,
         net712966, net712844, net712841, net712840, net712487, net712486,
         net712447, net712359, net783365, net780581, net762630, net760174,
         net758891, net755642, net755215, net753295, net749831, net749633,
         net749368, net746029, net742308, net740525, net738752, net736222,
         net732820, net732819, net731203, net727668, net720607, net717607,
         net717564, net714856, net714833, net714742, net714705, net714703,
         net714702, net714328, net714136, net713921, net713709, net750018,
         net727275, net718336, net717802, net717594, net715748, net715432,
         net715167, net714961, net714323, net714058, net713749, net713695,
         net786871, net755063, net749609, net742288, net742051, net720497,
         net720496, net715787, net715786, net715785, net715774, net715770,
         net715751, net715746, net812279, net812284, net812773, net812861,
         net812866, net812941, net812952, net812958, net826165, net713413,
         net712645, n18833, n18832, n18831, n18828, n18827, n18826, n18825,
         n18824, n18823, n18822, n18821, n18819, n18818, n18817, n18816,
         n18815, n18814, net839583, net780338, net717654, net713451, net713441,
         net712366, net780599, net780295, net780294, net716251, net712367,
         net873523, net804645, net795260, net780225, net765379, net760673,
         net760672, net755203, net740705, net729283, net729282, net727306,
         net714621, net714620, net714619, net714342, net714341, net714340,
         net714339, net714332, net714330, net714087, net714086, net714085,
         net714032, net714031, net714030, net713490, net713488, net713461,
         net713455, net713450, net713449, net713068, net713067, net713062,
         net712946, net712888, net712559, n18887, n18886, n18885, n18882,
         n18881, n18880, n18879, n18878, n18877, n18876, n18875, n18873,
         n18872, n18871, n18870, n18869, n18868, net795965, net795964,
         net762727, net755262, net752497, net750251, net750159, net737941,
         net727829, net727828, net727827, net718025, net717464, net715603,
         net715242, net715232, net714967, net714876, net714874, net714408,
         net714407, net714406, net714377, net714376, net714375, net714362,
         net714361, net714360, net714078, net713453, net712815, net712799,
         net712452, net742258, net741960, net741847, net739688, net724878,
         net724877, net718360, net718032, net717517, net717509, net717107,
         net713847, net713680, net812287, net804492, net750077, net749815,
         net749287, net745725, net745723, net742371, net742073, net740358,
         net740357, net740305, net740183, net739743, net739296, net720499,
         net720498, net718093, net718026, net717955, net715814, net715810,
         net715782, net715781, net715780, net715779, net715778, net715771,
         net715696, net715691, net715690, net715688, net715677, net715676,
         net715674, net715673, net715663, net715593, net715590, n22612, n22613,
         n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621,
         n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629,
         n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637,
         n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645,
         n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653,
         n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661,
         n22662, n22663, n22664, n22665, n22666, n22667, n22669, n22670,
         n22671, n22672, n22673, n22674, n22675, n22676, n22677, n22678,
         n22679, n22680, n22681, n22682, n22683, n22684, n22685, n22686,
         n22687, n22688, n22689, n22690, n22691, n22693, n22694, n22695,
         n22696, n22697, n22698, n22699, n22700, n22701, n22702, n22703,
         n22704, n22705, n22706, n22707, n22708, n22709, n22710, n22711,
         n22712, n22713, n22714, n22715, n22716, n22717, n22718, n22719,
         n22720, n22721, n22722, n22723, n22724, n22725, n22726, n22727,
         n22728, n22729, n22730, n22731, n22732, n22733, n22734, n22735,
         n22736, n22737, n22738, n22739, n22740, n22742, n22745, n22759,
         n22760, n22761, n22762, n22763, n22764, n22765, n22766, n22767,
         n22768, n22769, n22770, n22771, n22772, n22773, n22774, n22775,
         n22776, n22777, n22778, n22779, n22780, n22781, n22782, n22783,
         n22784, n22785, n22786, n22787, n22788, n22789, n22790, n22791,
         n22792, n22793, n22794, n22795, n22796, n22797, n22798, n22799,
         n22800, n22801, n22802, n22803, n22804, n22805, n22806, n22807,
         n22808, n22809, n22810, n22811, n22812, n22813, n22814, n22815,
         n22816, n22817, n22818, n22819, n22820, n22821, n22822, n22823,
         n22824, n22825, n22826, n22827, n22828, n22829, n22830, n22831,
         n22832, n22833, n22834, n22835, n22836, n22837, n22838, n22839,
         n22840, n22841, n22842, n22843, n22844, n22845, n22847, n22850,
         n22851, n22852, n22853, n22855, n22856, n22858, n22859, n22860,
         n22861, n22862, n22863, n22864, n22865, n22866, n22867, n22868,
         n22869, n22870, n22871, n22872, n22873, n22874, n22875, n22876,
         n22877, n22878, n22879, n22880, n22881, n22882, n22883, n22884,
         n22885, n22886, n22887, n22888, n22889, n22890, n22891, n22892,
         n22893, n22894, n22895, n22896, n22897, n22898, n22899, n22900,
         n22901, n22902, n22903, n22904, n22905, n22906, n22907, n22908,
         n22909, n22910, n22911, n22912, n22913, n22914, n22915, n22916,
         n22917, n22918, n22919, n22920, n22921, n22922, n22923, n22924,
         n22925, n22926, n22927, n22928, n22929, n22930, n22931, n22932,
         n22933, n22934, n22935, n22936, n22938, n22939, n22940, n22941,
         n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949,
         n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957,
         n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965,
         n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973,
         n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981,
         n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989,
         n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997,
         n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005,
         n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013,
         n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021,
         n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029,
         n23030, n23031, n23041, n23042, n23043, n23044, n23045, n23046,
         n23047, n23048, n23049, n23050, n23051, n23052, n23053, n23054,
         n23055, n23056, n23057, n23058, n23059, n23060, n23061, n23062,
         n23063, n23064, n23065, n23066, n23067, n23068, n23069, n23070,
         n23071, n23072, n23073, n23074, n23075, n23076, n23077, n23078,
         n23079, n23080, n23081, n23082, n23083, n23084, n23085, n23086,
         n23087, n23088, n23089, n23090, n23091, n23092, n23093, n23094,
         n23095, n23096, n23097, n23098, n23099, n23100, n23101, n23102,
         n23103, n23104, n23105, n23106, n23107, n23108, n23109, n23110,
         n23111, n23112, n23113, n23114, n23115, n23116, n23117, n23118,
         n23119, n23120, n23121, n23122, n23123, n23124, n23125, n23126,
         n23127, n23128, n23129, n23130, n23131, n23132, n23133, n23134,
         n23135, n23136, n23137, n23138, n23139, n23140, n23141, n23142,
         n23143, n23144, n23145, n23146, n23147, n23148, n23149, n23150,
         n23151, n23152, n23153, n23154, n23155, n23156, n23157, n23158,
         n23159, n23160, n23161, n23162, n23163, n23164, n23165, n23166,
         n23167, n23168, n23169, n23170, n23171, n23172, n23173, n23174,
         n23175, n23176, n23177, n23178, n23179, n23180, n23181, n23182,
         n23183, n23184, n23185, n23186, n23187, n23188, n23189, n23190,
         n23191, n23192, n23193, n23194, n23195, n23196, n23197, n23198,
         n23199, n23200, n23201, n23202, n23203, n23204, n23205, n23206,
         n23207, n23208, n23209, n23210, n23211, n23212, n23213, n23214,
         n23215, n23216, n23217, n23218, n23219, n23220, n23221, n23222,
         n23223, n23224, n23225, n23226, n23227, n23228, n23229, n23230,
         n23231, n23232, n23233, n23234, n23235, n23236, n23237, n23238,
         n23239, n23240, n23241, n23242, n23243, n23244, n23245, n23246,
         n23247, n23248, n23249, n23250, n23251, n23252, n23253, n23254,
         n23255, n23256, n23257, n23258, n23259, n23260, n23261, n23262,
         n23263, n23264, n23265, n23266, n23267, n23268, n23269, n23270,
         n23271, n23272, n23273, n23274, n23275, n23276, n23277, n23278,
         n23279, n23280, n23281, n23282, n23283, n23284, n23285, n23286,
         n23287, n23288, n23289, n23290, n23291, n23292, n23293, n23294,
         n23295, n23296, n23297, n23298, n23299, n23300, n23301, n23302,
         n23303, n23304, n23305, n23306, n23307, n23308, n23309, n23310,
         n23311, n23312, n23313, n23314, n23315, n23316, n23317, n23318,
         n23319, n23320, n23321, n23322, n23323, n23324, n23325, n23326,
         n23327, n23328, n23329, n23330, n23331, n23332, n23333, n23334,
         n23335, n23336, n23337, n23338, n23339, n23340, n23341, n23342,
         n23343, n23344, n23345, n23346, n23347, n23348, n23349, n23350,
         n23351, n23352, n23353, n23354, n23355, n23356, n23357, n23358,
         n23359, n23360, n23361, n23362, n23363, n23364, n23365, n23366,
         n23367, n23368, n23369, n23370, n23371, n23372, n23373, n23374,
         n23375, n23376, n23377, n23378, n23379, n23380, n23381, n23382,
         n23383, n23384, n23385, n23386, n23387, n23388, n23389, n23390,
         n23391, n23392, n23393, n23394, n23395, n23396, n23397, n23398,
         n23399, n23400, n23401, n23402, n23403, n23404, n23405, n23406,
         n23407, n23408, n23409, n23410, n23411, n23412, n23413, n23414,
         n23415, n23416, n23417, n23418, n23419, n23420, n23421, n23422,
         n23423, n23424, n23425, n23426, n23427, n23428, n23429, n23430,
         n23431, n23432, n23433, n23434, n23435, n23436, n23437, n23438,
         n23439, n23440, n23441, n23442, n23443, n23444, n23445, n23446,
         n23447, n23448, n23449, n23450, n23451, n23452, n23453, n23454,
         n23455, n23456, n23457, n23458, n23459, n23460, n23461, n23462,
         n23463, n23464, n23465, n23466, n23467, n23468, n23469, n23470,
         n23471, n23472, n23473, n23474, n23475, n23476, n23477, n23478,
         n23479, n23480, n23481, n23482, n23483, n23484, n23485, n23486,
         n23487, n23488, n23489, n23490, n23491, n23492, n23493, n23494,
         n23495, n23496, n23497, n23498, n23499, n23500, n23501, n23502,
         n23503, n23504, n23505, n23506, n23507, n23508, n23509, n23510,
         n23511, n23512, n23513, n23514, n23515, n23516, n23517, n23518,
         n23519, n23520, n23521, n23522, n23523, n23524, n23525, n23526,
         n23527, n23528, n23529, n23530, n23531, n23532, n23533, n23534,
         n23535, n23536, n23537, n23538, n23539, n23540, n23541, n23542,
         n23543, n23544, n23545, n23546, n23547, n23548, n23549, n23550,
         n23551, n23552, n23553, n23554, n23555, n23556, n23557, n23558,
         n23559, n23560, n23561, n23562, n23563, n23564, n23565, n23566,
         n23567, n23568, n23569, n23570, n23571, n23572, n23573, n23574,
         n23575, n23576, n23577, n23578, n23579, n23580, n23581, n23582,
         n23583, n23584, n23585, n23586, n23587, n23588, n23589, n23590,
         n23591, n23592, n23593, n23594, n23595, n23596, n23597, n23598,
         n23599, n23600, n23601, n23602, n23603, n23604, n23605, n23606,
         n23607, n23608, n23609, n23610, n23611, n23612, n23613, n23614,
         n23615, n23616, n23617, n23618, n23619, n23620, n23621, n23622,
         n23623, n23624, n23625, n23626, n23627, n23628, n23629, n23630,
         n23631, n23632, n23633, n23634, n23635, n23636, n23637, n23638,
         n23639, n23640, n23641, n23642, n23643, n23644, n23645, n23646,
         n23647, n23648, n23649, n23650, n23651, n23652, n23653, n23654,
         n23655, n23656, n23657, n23658, n23659, n23660, n23661, n23662,
         n23663, n23664, n23665, n23666, n23667, n23668, n23669, n23670,
         n23671, n23672, n23673, n23674, n23675, n23676, n23677, n23678,
         n23679, n23680, n23681, n23682, n23683, n23684, n23685, n23686,
         n23687, n23688, n23689, n23690, n23691, n23692, n23693, n23694,
         n23695, n23696, n23697, n23698, n23699, n23700, n23701, n23702,
         n23703, n23704, n23705, n23706, n23707, n23708, n23709, n23710,
         n23711, n23712, n23713, n23714, n23715, n23716, n23717, n23718,
         n23719, n23720, n23721, n23722, n23723, n23724, n23725, n23726,
         n23727, n23728, n23729, n23730, n23731, n23732, n23733, n23734,
         n23735, n23736, n23737, n23738, n23739, n23740, n23741, n23742,
         n23743, n23744, n23745, n23746, n23747, n23748, n23749, n23750,
         n23751, n23752, n23753, n23754, n23755, n23756, n23757, n23758,
         n23759, n23760, n23761, n23762, n23763, n23764, n23765, n23766,
         n23767, n23768, n23769, n23770, n23771, n23772, n23773, n23774,
         n23775, n23776, n23777, n23778, n23779, n23780, n23781, n23782,
         n23783, n23784, n23785, n23786, n23787, n23788, n23789, n23790,
         n23791, n23792, n23793, n23794, n23795, n23796, n23797, n23798,
         n23799, n23800, n23801, n23802, n23803, n23804, n23805, n23806,
         n23807, n23808, n23809, n23810, n23811, n23812, n23813, n23814,
         n23815, n23816, n23817, n23818, n23819, n23820, n23821, n23822,
         n23823, n23824, n23825, n23826, n23827, n23828, n23829, n23830,
         n23831, n23832, n23833, n23834, n23835, n23836, n23837, n23838,
         n23839, n23840, n23841, n23842, n23843, n23844, n23845, n23846,
         n23847, n23848, n23849, n23850, n23851, n23852, n23853, n23854,
         n23855, n23856, n23857, n23858, n23859, n23860, n23861, n23862,
         n23863, n23864, n23865, n23866, n23867, n23868, n23869, n23870,
         n23871, n23872, n23873, n23874, n23875, n23876, n23877, n23878,
         n23879, n23880, n23881, n23882, n23883, n23884, n23885, n23886,
         n23887, n23888, n23889, n23890, n23891, n23892, n23893, n23894,
         n23895, n23896, n23897, n23898, n23899, n23900, n23901, n23902,
         n23903, n23904, n23905, n23906, n23907, n23908, n23909, n23910,
         n23911, n23912, n23913, n23914, n23915, n23916, n23917, n23918,
         n23919, n23920, n23921, n23922, n23923, n23924, n23925, n23926,
         n23927, n23928, n23929, n23930, n23931, n23932, n23933, n23934,
         n23935, n23936, n23937, n23938, n23939, n23940, n23941, n23942,
         n23944, n23946, n23947, n23948, n23949, n23950, n23951, n23952,
         n23953, n23954, n23955, n23956, n23957, n23958, n23959, n23960,
         n23961, n23962, n23963, n23964, n23965, n23966, n23967, n23968,
         n23969, n23970, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24102, n24103, n24104, n24105, n24106, n24107,
         n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
         n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123,
         n24124, n24125, n24126, n24128, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24175, n24176, n24177, n24178,
         n24179, n24190, n24191, n24192, n24193, n24194, n24195, n24196,
         n24197, n24198, n24199, n24200, n24201, n24202, n24203, n24204,
         n24205, n24206, n24209, n24210, n24211, n24212, n24213, n24214,
         n24215, n24216, n24217, n24218, n24219, n24220, n24221, n24222,
         n24223, n24224, n24225, n24226, n24227, n24228, n24229, n24230,
         n24231, n24232, n24233, n24234, n24235, n24236, n24237, n24238,
         n24239, n24240, n24241, n24242, n24243, n24244, n24245, n24246,
         n24247, n24248, n24249, n24250, n24251, n24252, n24253, n24254,
         n24255, n24256, n24257, n24258, n24259, n24260, n24261, n24262,
         n24263, n24264, n24265, n24266, n24267, n24268, n24269, n24270,
         n24271, n24272, n24273, n24274, n24275, n24276, n24277, n24278,
         n24279, n24280, n24281, n24282, n24283, n24284, n24285, n24286,
         n24287, n24288, n24289, n24290, n24291, n24292, n24293, n24294,
         n24295, n24296, n24297, n24298, n24299, n24300, n24301, n24302,
         n24303, n24304, n24305, n24306, n24307, n24308, n24309, n24310,
         n24311, n24312, n24313, n24314, n24315, n24316, n24317, n24318,
         n24319, n24320, n24321, n24322, n24323, n24324, n24325, n24326,
         n24327, n24328, n24329, n24330, n24331, n24332, n24333, n24334,
         n24335, n24336, n24337, n24338, n24339, n24340, n24341, n24342,
         n24343, n24344, n24345, n24346, n24347, n24348, n24349, n24350,
         n24351, n24352, n24353, n24354, n24355, n24356, n24357, n24358,
         n24359, n24360, n24361, n24362, n24363, n24364, n24365, n24366,
         n24367, n24368, n24369, n24370, n24371, n24372, n24373, n24374,
         n24375, n24376, n24377, n24378, n24379, n24380, n24381, n24382,
         n24383, n24384, n24385, n24386, n24387, n24388, n24389, n24390,
         n24391, n24392, n24393, n24394, n24395, n24396, n24397, n24398,
         n24399, n24400, n24401, n24402, n24403, n24404, n24405, n24406,
         n24407, n24408, n24409, n24410, n24411, n24412, n24413, n24414,
         n24415, n24416, n24417, n24418, n24419, n24420, n24421, n24422,
         n24423, n24424, n24425, n24426, n24427, n24428, n24429, n24430,
         n24431, n24432, n24433, n24434, n24435, n24436, n24437, n24438,
         n24439, n24440, n24441, n24442, n24443, n24444, n24445, n24446,
         n24447, n24448, n24449, n24450, n24451, n24452, n24453, n24454,
         n24455, n24456, n24457, n24458, n24459, n24460, n24461, n24462,
         n24463, n24464, n24465, n24466, n24467, n24468, n24469, n24470,
         n24471, n24472, n24473, n24474, n24475, n24476, n24477, n24478,
         n24479, n24480, n24481, n24482, n24483, n24484, n24485, n24486,
         n24487, n24488, n24489, n24490, n24491, n24492, n24493, n24494,
         n24495, n24496, n24497, n24498, n24499, n24500, n24501, n24502,
         n24503, n24504, n24505, n24506, n24507, n24508, n24509, n24510,
         n24511, n24512, n24513, n24514, n24515, n24516, n24517, n24518,
         n24519, n24520, n24521, n24522, n24523, n24524, n24525, n24526,
         n24527, n24528, n24529, n24530, n24531, n24532, n24533, n24534,
         n24535, n24536, n24537, n24538, n24539, n24540, n24541, n24542,
         n24543, n24544, n24545, n24546, n24547, n24548, n24549, n24550,
         n24551, n24552, n24553, n24554, n24555, n24556, n24557, n24558,
         n24559, n24560, n24561, n24562, n24563, n24564, n24565, n24566,
         n24567, n24568, n24569, n24570, n24571, n24572, n24573, n24574,
         n24575, n24576, n24577, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785;
  wire   [1:0] s_MEM_LOAD_TYPE;
  wire   [1:0] s_WB_MUX_CONTROL;
  wire   [31:0] s_IFID_IR;
  wire   [31:0] s_MEMWB_IR;
  wire   [31:0] \core_inst/ps_EXMEM_DATA_IN ;
  wire   [31:0] \core_inst/s_IF_OUT_IR_OUT ;
  wire  
         [31:0] \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p 
;
  tri   [31:0] DRAM_INTERFACE;
  tri   \core_inst/s_DRAM_DLX_OUT[16] ;
  tri   \core_inst/s_DRAM_DLX_OUT[17] ;
  tri   \core_inst/s_DRAM_DLX_OUT[18] ;
  tri   \core_inst/s_DRAM_DLX_OUT[19] ;
  tri   \core_inst/s_DRAM_DLX_OUT[20] ;
  tri   \core_inst/s_DRAM_DLX_OUT[21] ;
  tri   \core_inst/s_DRAM_DLX_OUT[22] ;
  tri   \core_inst/s_DRAM_DLX_OUT[23] ;
  tri   \core_inst/s_DRAM_DLX_OUT[24] ;
  tri   \core_inst/s_DRAM_DLX_OUT[25] ;
  tri   \core_inst/s_DRAM_DLX_OUT[26] ;
  tri   \core_inst/s_DRAM_DLX_OUT[27] ;
  tri   \core_inst/s_DRAM_DLX_OUT[28] ;
  tri   \core_inst/s_DRAM_DLX_OUT[29] ;
  tri   \core_inst/s_DRAM_DLX_OUT[30] ;
  tri   \core_inst/s_DRAM_DLX_OUT[31] ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_0/s_top ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_1/s_top ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_2/s_top ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_3/s_top ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_4/s_top ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_5/s_top ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_6/s_top ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_7/s_top ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_8/s_top ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_9/s_top ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_10/s_top ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_11/s_top ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_12/s_top ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_13/s_top ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_14/s_top ;
  tri   \core_inst/MEM/MUX_LOAD/MUX_BIT_15/s_top ;
  assign \core_inst/s_IF_OUT_IR_OUT  [0] = ROM_INTERFACE[0];
  assign \core_inst/s_IF_OUT_IR_OUT  [1] = ROM_INTERFACE[1];
  assign \core_inst/s_IF_OUT_IR_OUT  [2] = ROM_INTERFACE[2];
  assign \core_inst/s_IF_OUT_IR_OUT  [3] = ROM_INTERFACE[3];
  assign \core_inst/s_IF_OUT_IR_OUT  [4] = ROM_INTERFACE[4];
  assign \core_inst/s_IF_OUT_IR_OUT  [5] = ROM_INTERFACE[5];
  assign \core_inst/s_IF_OUT_IR_OUT  [6] = ROM_INTERFACE[6];
  assign \core_inst/s_IF_OUT_IR_OUT  [7] = ROM_INTERFACE[7];
  assign \core_inst/s_IF_OUT_IR_OUT  [8] = ROM_INTERFACE[8];
  assign \core_inst/s_IF_OUT_IR_OUT  [9] = ROM_INTERFACE[9];
  assign \core_inst/s_IF_OUT_IR_OUT  [10] = ROM_INTERFACE[10];
  assign \core_inst/s_IF_OUT_IR_OUT  [11] = ROM_INTERFACE[11];
  assign \core_inst/s_IF_OUT_IR_OUT  [12] = ROM_INTERFACE[12];
  assign \core_inst/s_IF_OUT_IR_OUT  [13] = ROM_INTERFACE[13];
  assign \core_inst/s_IF_OUT_IR_OUT  [14] = ROM_INTERFACE[14];
  assign \core_inst/s_IF_OUT_IR_OUT  [15] = ROM_INTERFACE[15];
  assign \core_inst/s_IF_OUT_IR_OUT  [16] = ROM_INTERFACE[16];
  assign \core_inst/s_IF_OUT_IR_OUT  [17] = ROM_INTERFACE[17];
  assign \core_inst/s_IF_OUT_IR_OUT  [18] = ROM_INTERFACE[18];
  assign \core_inst/s_IF_OUT_IR_OUT  [19] = ROM_INTERFACE[19];
  assign \core_inst/s_IF_OUT_IR_OUT  [20] = ROM_INTERFACE[20];
  assign \core_inst/s_IF_OUT_IR_OUT  [21] = ROM_INTERFACE[21];
  assign \core_inst/s_IF_OUT_IR_OUT  [22] = ROM_INTERFACE[22];
  assign \core_inst/s_IF_OUT_IR_OUT  [23] = ROM_INTERFACE[23];
  assign \core_inst/s_IF_OUT_IR_OUT  [24] = ROM_INTERFACE[24];
  assign \core_inst/s_IF_OUT_IR_OUT  [25] = ROM_INTERFACE[25];
  assign \core_inst/s_IF_OUT_IR_OUT  [26] = ROM_INTERFACE[26];
  assign \core_inst/s_IF_OUT_IR_OUT  [27] = ROM_INTERFACE[27];
  assign \core_inst/s_IF_OUT_IR_OUT  [28] = ROM_INTERFACE[28];
  assign \core_inst/s_IF_OUT_IR_OUT  [29] = ROM_INTERFACE[29];
  assign \core_inst/s_IF_OUT_IR_OUT  [30] = ROM_INTERFACE[30];
  assign \core_inst/s_IF_OUT_IR_OUT  [31] = ROM_INTERFACE[31];
  assign ROM_ADDRESS[3] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_up_network_p[1] ;
  assign ROM_ADDRESS[2] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_g[2] ;
  assign ROM_ADDRESS[1] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [1];
  assign ROM_ADDRESS[4] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [4];
  assign ROM_ADDRESS[5] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [5];
  assign ROM_ADDRESS[6] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [6];
  assign ROM_ADDRESS[7] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [7];
  assign ROM_ADDRESS[8] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [8];
  assign ROM_ADDRESS[9] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [9];
  assign ROM_ADDRESS[10] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [10];
  assign ROM_ADDRESS[11] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [11];
  assign ROM_ADDRESS[12] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [12];
  assign ROM_ADDRESS[13] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [13];
  assign ROM_ADDRESS[14] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [14];
  assign ROM_ADDRESS[15] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [15];
  assign ROM_ADDRESS[16] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [16];
  assign ROM_ADDRESS[17] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [17];
  assign ROM_ADDRESS[18] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [18];
  assign ROM_ADDRESS[19] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [19];
  assign ROM_ADDRESS[20] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [20];
  assign ROM_ADDRESS[21] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [21];
  assign ROM_ADDRESS[22] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [22];
  assign ROM_ADDRESS[23] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [23];
  assign ROM_ADDRESS[24] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [24];
  assign ROM_ADDRESS[25] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [25];
  assign ROM_ADDRESS[26] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [26];
  assign ROM_ADDRESS[27] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [27];
  assign ROM_ADDRESS[28] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [28];
  assign ROM_ADDRESS[29] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p  [29];
  assign ROM_ADDRESS[0] = \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/CLA_PG_NET/N1 ;
  assign ROM_ADDRESS[31] = \core_inst/IF_stage/PLUS4_ADDER/RES_GENERATOR/CSA_15/sum_rca_0[1] ;
  assign ROM_ADDRESS[30] = \core_inst/IF_stage/PLUS4_ADDER/RES_GENERATOR/CSA_15/RCA_1/cout_tmp[0] ;
  assign DRAM_ADDRESS[0] = \core_inst/MEMWB_ALUOUT/DFF_0/N3 ;
  assign DRAM_ADDRESS[1] = \core_inst/MEMWB_ALUOUT/DFF_1/N3 ;
  assign DRAM_ADDRESS[2] = \core_inst/MEMWB_ALUOUT/DFF_2/N3 ;
  assign DRAM_ADDRESS[3] = \core_inst/MEMWB_ALUOUT/DFF_3/N3 ;
  assign DRAM_ADDRESS[4] = \core_inst/MEMWB_ALUOUT/DFF_4/N3 ;
  assign DRAM_ADDRESS[5] = \core_inst/MEMWB_ALUOUT/DFF_5/N3 ;
  assign DRAM_ADDRESS[6] = \core_inst/MEMWB_ALUOUT/DFF_6/N3 ;
  assign DRAM_ADDRESS[7] = \core_inst/MEMWB_ALUOUT/DFF_7/N3 ;
  assign DRAM_ADDRESS[8] = \core_inst/MEMWB_ALUOUT/DFF_8/N3 ;
  assign DRAM_ADDRESS[9] = \core_inst/MEMWB_ALUOUT/DFF_9/N3 ;
  assign DRAM_ADDRESS[10] = \core_inst/MEMWB_ALUOUT/DFF_10/N3 ;
  assign DRAM_ADDRESS[11] = \core_inst/MEMWB_ALUOUT/DFF_11/N3 ;
  assign DRAM_ADDRESS[12] = \core_inst/MEMWB_ALUOUT/DFF_12/N3 ;
  assign DRAM_ADDRESS[13] = \core_inst/MEMWB_ALUOUT/DFF_13/N3 ;
  assign DRAM_ADDRESS[14] = \core_inst/MEMWB_ALUOUT/DFF_14/N3 ;
  assign DRAM_ADDRESS[15] = \core_inst/MEMWB_ALUOUT/DFF_15/N3 ;
  assign DRAM_ADDRESS[16] = \core_inst/MEMWB_ALUOUT/DFF_16/N3 ;
  assign DRAM_ADDRESS[17] = \core_inst/MEMWB_ALUOUT/DFF_17/N3 ;
  assign DRAM_ADDRESS[18] = \core_inst/MEMWB_ALUOUT/DFF_18/N3 ;
  assign DRAM_ADDRESS[19] = \core_inst/MEMWB_ALUOUT/DFF_19/N3 ;
  assign DRAM_ADDRESS[20] = \core_inst/MEMWB_ALUOUT/DFF_20/N3 ;
  assign DRAM_ADDRESS[21] = \core_inst/MEMWB_ALUOUT/DFF_21/N3 ;
  assign DRAM_ADDRESS[22] = \core_inst/MEMWB_ALUOUT/DFF_22/N3 ;
  assign DRAM_ADDRESS[23] = \core_inst/MEMWB_ALUOUT/DFF_23/N3 ;
  assign DRAM_ADDRESS[24] = \core_inst/MEMWB_ALUOUT/DFF_24/N3 ;
  assign DRAM_ADDRESS[25] = \core_inst/MEMWB_ALUOUT/DFF_25/N3 ;
  assign DRAM_ADDRESS[26] = \core_inst/MEMWB_ALUOUT/DFF_26/N3 ;
  assign DRAM_ADDRESS[27] = \core_inst/MEMWB_ALUOUT/DFF_27/N3 ;
  assign DRAM_ADDRESS[28] = \core_inst/MEMWB_ALUOUT/DFF_28/N3 ;
  assign DRAM_ADDRESS[29] = \core_inst/MEMWB_ALUOUT/DFF_29/N3 ;
  assign DRAM_ADDRESS[30] = \core_inst/MEMWB_ALUOUT/DFF_30/N3 ;
  assign DRAM_ADDRESS[31] = \core_inst/MEMWB_ALUOUT/DFF_31/N3 ;
  assign ROM_EN = 1'b1;
  assign DRAM_EN = 1'b1;
  assign DRAM_READNOTWRITE = \core_inst/N65 ;

  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n1755) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_31/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_31/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net741582), .QN(n4347) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_31/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_31/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24773), .QN(n4346) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_0/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_0/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24781), .QN(n4421) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_10/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_10/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24806), .QN(n4415) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_11/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_11/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24607), .QN(n4412) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_12/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_12/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net740710), .QN(n4409) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_27/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_27/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24783), .QN(n4361) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_17/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_17/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n25317), .QN(n4394) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_25/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_25/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24603), .QN(n4367) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_22/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_22/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n5664), .QN(n25282) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_30/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_30/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_30/N3 ), .QN(n1734) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_30/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_30/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n25328) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_14/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_14/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_14/N3 ), .QN(n1732) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_14/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_14/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n25327) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_29/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_29/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24604), .QN(n4355) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_26/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_26/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_26/N3 ), .QN(n1728) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_26/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_26/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24605), .QN(n4364) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_8/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_8/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net741580), .QN(n4331) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_23/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_23/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_23/N3 ), .QN(n1724) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_23/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_23/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n25318), .QN(n4373) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_18/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_18/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n25330), .QN(n4391) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_24/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_24/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n25337) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_19/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_19/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net741301), .QN(n4388) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_28/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_28/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24784), .QN(n4358) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_9/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_9/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24809), .QN(n4325) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_13/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_13/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_13/N3 ), .QN(n1712) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_13/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_13/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24782), .QN(n4406) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_15/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_15/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24606), .QN(n4400) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_16/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_16/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24807), .QN(n4397) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_6/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_6/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_6/N3 ), .QN(n1706) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_6/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_6/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24780), .QN(n4337) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_4/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_4/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24602), .QN(n4343) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_20/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_20/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24808), .QN(n4382) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_2/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_2/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_2/N3 ), .QN(n1700) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_2/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_2/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net741464), .QN(n4385) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_21/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_21/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n25329), .QN(n4379) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_7/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_7/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net365821), .QN(n24609) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_5/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_5/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net365826), .QN(n25339) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_3/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net741329), .QN(n4352) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_1/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_1/N3 ), .QN(n1690) );
  DFFR_X1 \core_inst/MEMWB_ALUOUT/DFF_1/data_reg  ( .D(
        \core_inst/MEMWB_ALUOUT/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n25319), .QN(n4418) );
  DFFR_X1 \core_inst/IFID_IR/DFF_9/data_reg  ( .D(\core_inst/IFID_IR/DFF_9/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n18066) );
  DFFR_X1 \core_inst/IFID_IR/DFF_8/data_reg  ( .D(\core_inst/IFID_IR/DFF_8/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n18065) );
  DFFR_X1 \core_inst/IFID_IR/DFF_7/data_reg  ( .D(\core_inst/IFID_IR/DFF_7/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n18064) );
  DFFR_X1 \core_inst/IFID_IR/DFF_6/data_reg  ( .D(\core_inst/IFID_IR/DFF_6/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n18063) );
  DFFR_X1 \core_inst/IFID_IR/DFF_5/data_reg  ( .D(\core_inst/IFID_IR/DFF_5/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n18062), .QN(n24677) );
  DFFR_X1 \core_inst/IFID_IR/DFF_4/data_reg  ( .D(\core_inst/IFID_IR/DFF_4/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n14210), .QN(n24785) );
  DFFR_X1 \core_inst/IFID_IR/DFF_31/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_31/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n14191), 
        .QN(n24612) );
  DFFR_X1 \core_inst/IFID_IR/DFF_21/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_21/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_IFID_IR[21]), .QN(net741353) );
  DFFR_X1 \core_inst/IFID_IR/DFF_17/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_17/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_IFID_IR[17]), .QN(net741620) );
  DFFR_X1 \core_inst/IFID_IR/DFF_15/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_15/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n25588), 
        .QN(n1684) );
  DFFR_X1 \core_inst/IFID_IR/DFF_12/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_12/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(n13165) );
  DFFR_X1 \core_inst/IFID_IR/DFF_11/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_11/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n25335)
         );
  DFFR_X1 \core_inst/IFID_IR/DFF_10/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_10/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        net873523) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_9/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_9/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n1678) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_8/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_8/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n1677) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_24/data_reg  ( .D(n22702), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net366410), .QN(net718069) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_23/data_reg  ( .D(n22867), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net342961), .QN(net718070) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_22/data_reg  ( .D(n22801), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net342954), .QN(net718006) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_21/data_reg  ( .D(net712344), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(net342963), .QN(n25589) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_20/data_reg  ( .D(n22945), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net342852), .QN(net717830) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_18/data_reg  ( .D(n22703), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net342960), .QN(net717952) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_15/data_reg  ( .D(n22939), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18058) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_15/data_reg  ( .D(n22939), .CK(DLX_CLK), 
        .RN(DLX_RST), .QN(n25358) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_14/data_reg  ( .D(n26743), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18056) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_13/data_reg  ( .D(n26742), .CK(DLX_CLK), 
        .RN(DLX_RST), .QN(n1659) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_12/data_reg  ( .D(net712313), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n18055) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_11/data_reg  ( .D(n26741), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18054) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_11/data_reg  ( .D(n26741), .CK(DLX_CLK), 
        .RN(DLX_RST), .QN(n1655) );
  DFFR_X1 \core_inst/MEMWB_IR/DFF_20/data_reg  ( .D(
        \core_inst/MEMWB_IR/DFF_20/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n25593) );
  DFFR_X1 \core_inst/EXMEM_IR/DFF_19/data_reg  ( .D(
        \core_inst/EXMEM_IR/DFF_19/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_IR/DFF_19/N3 ), .QN(n1651) );
  DFFR_X1 \core_inst/MEMWB_IR/DFF_19/data_reg  ( .D(
        \core_inst/MEMWB_IR/DFF_19/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_MEMWB_IR[19]), .QN(n25582) );
  DFFR_X1 \core_inst/EXMEM_IR/DFF_18/data_reg  ( .D(
        \core_inst/EXMEM_IR/DFF_18/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n18053), .QN(n1649) );
  DFFR_X1 \core_inst/MEMWB_IR/DFF_17/data_reg  ( .D(
        \core_inst/MEMWB_IR/DFF_17/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n24336), .QN(n25584) );
  DFFR_X1 \core_inst/MEMWB_IR/DFF_16/data_reg  ( .D(
        \core_inst/MEMWB_IR/DFF_16/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n24315), .QN(n25583) );
  DFFR_X1 \core_inst/EXMEM_IR/DFF_15/data_reg  ( .D(
        \core_inst/EXMEM_IR/DFF_15/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_IR/DFF_15/N3 ), .QN(n1643) );
  DFFR_X1 \core_inst/MEMWB_IR/DFF_15/data_reg  ( .D(
        \core_inst/MEMWB_IR/DFF_15/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_MEMWB_IR[15]), .QN(net749230) );
  DFFR_X1 \core_inst/EXMEM_IR/DFF_14/data_reg  ( .D(
        \core_inst/EXMEM_IR/DFF_14/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_IR/DFF_14/N3 ), .QN(n1641) );
  DFFR_X1 \core_inst/MEMWB_IR/DFF_14/data_reg  ( .D(
        \core_inst/MEMWB_IR/DFF_14/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_MEMWB_IR[14]) );
  DFFR_X1 \core_inst/MEMWB_IR/DFF_13/data_reg  ( .D(
        \core_inst/MEMWB_IR/DFF_13/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_MEMWB_IR[13]) );
  DFFR_X1 \core_inst/MEMWB_IR/DFF_12/data_reg  ( .D(
        \core_inst/MEMWB_IR/DFF_12/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_MEMWB_IR[12]) );
  DFFR_X1 \core_inst/MEMWB_IR/DFF_11/data_reg  ( .D(
        \core_inst/MEMWB_IR/DFF_11/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_MEMWB_IR[11]), .QN(net749551) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_0/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_0/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n18052) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_1/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n18051) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_2/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_2/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n18050) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_3/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        net741306) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_4/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_4/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n24815) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_5/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_5/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n1628) );
  DFFR_X1 \core_inst/EXMEM_IR/DFF_29/data_reg  ( .D(
        \core_inst/EXMEM_IR/DFF_29/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net334510), .QN(net742046) );
  DFFR_X1 \core_inst/MEMWB_IR/DFF_29/data_reg  ( .D(net742047), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(s_MEMWB_IR[29]), .QN(net718098) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_31/data_reg  ( .D(
        \core_inst/IDEX_IR/DFF_31/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net741345), .QN(n14382) );
  DFFR_X1 \core_inst/MEMWB_IR/DFF_31/data_reg  ( .D(net89524), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n18047) );
  DFFR_X1 \cu_inst/EX/DFF_0/data_reg  ( .D(net710357), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(\cu_inst/MEM/DFF_0/N3 ) );
  DFFR_X1 \cu_inst/MEM/DFF_0/data_reg  ( .D(\cu_inst/MEM/DFF_0/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(\cu_inst/WB/DFF_0/N3 ) );
  DFFR_X1 \cu_inst/WB/DFF_0/data_reg  ( .D(\cu_inst/WB/DFF_0/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n18046) );
  DFFR_X1 \core_inst/MEMWB_IR/DFF_28/data_reg  ( .D(n25581), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(s_MEMWB_IR[28]), .QN(net718138) );
  DFFR_X1 \cu_inst/EX/DFF_18/data_reg  ( .D(\cu_inst/EX/DFF_18/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(s_EX_BRANCH_TYPE) );
  DFFR_X1 \cu_inst/EX/DFF_2/data_reg  ( .D(net710357), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(\cu_inst/MEM/DFF_2/N3 ) );
  DFFR_X1 \cu_inst/MEM/DFF_2/data_reg  ( .D(\cu_inst/MEM/DFF_2/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(\cu_inst/WB/DFF_2/N3 ) );
  DFFR_X1 \cu_inst/WB/DFF_2/data_reg  ( .D(\cu_inst/WB/DFF_2/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(s_WB_MUX_CONTROL[1]), .QN(n24679) );
  DFFR_X1 \cu_inst/EX/DFF_9/data_reg  ( .D(\cu_inst/EX/DFF_9/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(s_EX_IS_BRANCH), .QN(net740645) );
  DFFR_X1 \core_inst/EXMEM_IR/DFF_30/data_reg  ( .D(
        \core_inst/EXMEM_IR/DFF_30/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_IR/DFF_30/N3 ), .QN(\cu_inst/FW_UNIT/ITD_EXMEM/N14 )
         );
  DFFR_X1 \core_inst/MEMWB_IR/DFF_30/data_reg  ( .D(
        \core_inst/MEMWB_IR/DFF_30/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_MEMWB_IR[30]), .QN(net718111) );
  DFFR_X1 \cu_inst/EX/DFF_6/data_reg  ( .D(\cu_inst/EX/DFF_6/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(\cu_inst/MEM/DFF_6/N3 ) );
  DFFR_X1 \cu_inst/MEM/DFF_6/data_reg  ( .D(\cu_inst/MEM/DFF_6/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(s_MEM_SIGNED_LOAD) );
  DFFR_X1 \cu_inst/EX/DFF_5/data_reg  ( .D(\cu_inst/EX/DFF_5/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(\cu_inst/MEM/DFF_5/N3 ) );
  DFFR_X1 \cu_inst/MEM/DFF_5/data_reg  ( .D(\cu_inst/MEM/DFF_5/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(s_MEM_LOAD_TYPE[1]) );
  DFFR_X1 \cu_inst/EX/DFF_4/data_reg  ( .D(\cu_inst/EX/DFF_4/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(\cu_inst/MEM/DFF_4/N3 ) );
  DFFR_X1 \cu_inst/MEM/DFF_4/data_reg  ( .D(\cu_inst/MEM/DFF_4/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(s_MEM_LOAD_TYPE[0]), .QN(n24774) );
  DFFR_X1 \cu_inst/EX/DFF_7/data_reg  ( .D(\cu_inst/EX/DFF_7/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(n1600) );
  DFFR_X1 \cu_inst/EX/DFF_3/data_reg  ( .D(\cu_inst/EX/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(\cu_inst/MEM/DFF_3/N3 ) );
  DFFR_X1 \cu_inst/MEM/DFF_3/data_reg  ( .D(\cu_inst/MEM/DFF_3/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(\cu_inst/WB/DFF_3/N3 ) );
  DFFR_X1 \cu_inst/EX/DFF_1/data_reg  ( .D(\cu_inst/EX/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(\cu_inst/MEM/DFF_1/N3 ) );
  DFFR_X1 \cu_inst/MEM/DFF_1/data_reg  ( .D(\cu_inst/MEM/DFF_1/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(\cu_inst/WB/DFF_1/N3 ) );
  DFFR_X1 \cu_inst/WB/DFF_1/data_reg  ( .D(\cu_inst/WB/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(s_WB_MUX_CONTROL[0]), .QN(n24678) );
  DFFR_X1 \core_inst/EXMEM_RF_ADDR_DEST/DFF_4/data_reg  ( .D(
        \core_inst/EXMEM_RF_ADDR_DEST/DFF_4/N3 ), .CK(DLX_CLK), .RN(DLX_RST), 
        .Q(\core_inst/MEMWB_RF_ADDR_DEST/DFF_4/N3 ) );
  DFFR_X1 \core_inst/MEMWB_RF_ADDR_DEST/DFF_4/data_reg  ( .D(
        \core_inst/MEMWB_RF_ADDR_DEST/DFF_4/N3 ), .CK(DLX_CLK), .RN(DLX_RST), 
        .Q(n18042) );
  DFFR_X1 \core_inst/MEMWB_RF_ADDR_DEST/DFF_3/data_reg  ( .D(
        \core_inst/MEMWB_RF_ADDR_DEST/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), 
        .Q(n18041) );
  DFFR_X1 \core_inst/EXMEM_RF_ADDR_DEST/DFF_2/data_reg  ( .D(
        \core_inst/EXMEM_RF_ADDR_DEST/DFF_2/N3 ), .CK(DLX_CLK), .RN(DLX_RST), 
        .Q(\core_inst/MEMWB_RF_ADDR_DEST/DFF_2/N3 ) );
  DFFR_X1 \core_inst/MEMWB_RF_ADDR_DEST/DFF_2/data_reg  ( .D(
        \core_inst/MEMWB_RF_ADDR_DEST/DFF_2/N3 ), .CK(DLX_CLK), .RN(DLX_RST), 
        .Q(n18040) );
  DFFR_X1 \core_inst/EXMEM_RF_ADDR_DEST/DFF_1/data_reg  ( .D(
        \core_inst/EXMEM_RF_ADDR_DEST/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), 
        .Q(\core_inst/MEMWB_RF_ADDR_DEST/DFF_1/N3 ) );
  DFFR_X1 \core_inst/MEMWB_RF_ADDR_DEST/DFF_1/data_reg  ( .D(
        \core_inst/MEMWB_RF_ADDR_DEST/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), 
        .Q(n18039) );
  DFFR_X1 \core_inst/EXMEM_RF_ADDR_DEST/DFF_0/data_reg  ( .D(
        \core_inst/EXMEM_RF_ADDR_DEST/DFF_0/N3 ), .CK(DLX_CLK), .RN(DLX_RST), 
        .Q(\core_inst/MEMWB_RF_ADDR_DEST/DFF_0/N3 ) );
  DFFR_X1 \core_inst/MEMWB_RF_ADDR_DEST/DFF_0/data_reg  ( .D(
        \core_inst/MEMWB_RF_ADDR_DEST/DFF_0/N3 ), .CK(DLX_CLK), .RN(DLX_RST), 
        .Q(n18038) );
  DFFR_X1 \cu_inst/EX/DFF_12/data_reg  ( .D(\cu_inst/EX/DFF_12/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(net741603) );
  DFFR_X1 \cu_inst/EX/DFF_13/data_reg  ( .D(\cu_inst/EX/DFF_13/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(net741531) );
  DFFR_X1 \cu_inst/EX/DFF_14/data_reg  ( .D(\cu_inst/EX/DFF_14/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(net741282), .QN(net366211) );
  DFFR_X1 \cu_inst/EX/DFF_15/data_reg  ( .D(\cu_inst/EX/DFF_15/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(net741307), .QN(net366479) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_0/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_0/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_0/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_0/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_0/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n18036) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18035), .QN(n24999) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18034), .QN(n25250) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18033), .QN(n25201) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18032), .QN(n24971) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18031), .QN(n25175) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24627) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24628) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18028), .QN(n25153) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18027), .QN(n25145) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18026), .QN(n25107) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18025), .QN(n24892) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18024), .QN(n25263) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18023), .QN(n25098) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18022), .QN(n25271) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18021), .QN(n24850) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3131) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3124) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3125) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3117) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3107) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3118) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3102) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3103) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24695), .QN(n3097) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3098) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3108) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24686), .QN(n3090) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24697), .QN(n3134) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24696), .QN(n3135) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3130) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_0/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3089) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_0/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_0/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [0]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_0/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_0/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24587), .QN(n4422) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_1/data_reg  ( .D(net812866), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n18020) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_1/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_1/N3 ) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_1/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_1/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_1/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n18019) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18018), .QN(n25000) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18017), .QN(n25251) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18016), .QN(n25202) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18015), .QN(n24972) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18014), .QN(n25176) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24629) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24630) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18011), .QN(n25154) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18010), .QN(n25146) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18009), .QN(n25108) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18008), .QN(n24893) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18007), .QN(n25264) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18006), .QN(n25099) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18005), .QN(n25272) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18004), .QN(n24851) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2716) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2712) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2713) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2709) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2702) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2710) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2699) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2700) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24698), .QN(n2696) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2697) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2703) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24687), .QN(n2694) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24700), .QN(n2718) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24699), .QN(n2719) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2715) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_1/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2693) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_1/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [1]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_1/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net366126) );
  DFFR_X1 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_2/data_reg  ( .D(
        \core_inst/IF_stage/PROGRAM_COUNTER/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_g[2] ), .QN(n1498) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_2/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_2/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_2/N3 ) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_2/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_2/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_2/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_2/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_2/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n18003) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24674) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18001), .QN(n25314) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n18000), .QN(n25304) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17999), .QN(n24978) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17998), .QN(n25286) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24623) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24675) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17995), .QN(n24951) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24594) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24676) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17992), .QN(n24903) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24737), .QN(n1481) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17991), .QN(n25306) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17990), .QN(n25313) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17989), .QN(n25284) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2320) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2316) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2317) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2313) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2306) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2314) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2303) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2304) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2300) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2301) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24736), .QN(n2307) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2298) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2322) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24596), .QN(n2323) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2319) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_2/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_2/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2297) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_2/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_2/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [2]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_2/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_2/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n5707), .QN(net740649) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_3/data_reg  ( .D(
        \core_inst/IFID_NPC/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n17988)
         );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_3/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_3/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_3/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n17987) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24649) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17985), .QN(n25257) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17984), .QN(n25047) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17983), .QN(n24979) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17982), .QN(n25182) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24651) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24650) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17979), .QN(n25040) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24652) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24588) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17976), .QN(n24912) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24805), .QN(n1442) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17975), .QN(n24889) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17974), .QN(n24844) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17973), .QN(n25036) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2212) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2208) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2209) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2205) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24791), .QN(n2198) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2206) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2195) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2196) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2192) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2193) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24599), .QN(n2199) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2190) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2214) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24725), .QN(n2215) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2211) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_3/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_3/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2189) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_3/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [3]) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_4/data_reg  ( .D(n23981), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n22698) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_4/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_4/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_4/N3 ) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_4/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_4/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_4/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_4/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_4/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n17971) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17970), .QN(n25019) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17969), .QN(n25045) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17968), .QN(n24777) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17967), .QN(n25044) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17966), .QN(n25080) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17965), .QN(n24775) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17964), .QN(n24776) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17963), .QN(n25041) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n14393), .QN(n25152) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17962), .QN(n25128) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17961), .QN(n24915) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n25326) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17960), .QN(n25039) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17959), .QN(n25281) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17958), .QN(n24857) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24804), .QN(n2176) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2172) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2173) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2169) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2162) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2170) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2159) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2160) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24789), .QN(n2156) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2157) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2163) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24788), .QN(n2154) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24728), .QN(n2178) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24727), .QN(n2179) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24793), .QN(n2175) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_4/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_4/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2153) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_4/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_4/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17957) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_4/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_4/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [4]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_4/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_4/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net741305), .QN(n4344) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_5/data_reg  ( .D(
        \core_inst/IFID_NPC/DFF_5/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n17956)
         );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_5/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_5/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_5/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_5/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_5/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n17955) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24668) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17953), .QN(n25288) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17952), .QN(n25277) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17951), .QN(n24980) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17950), .QN(n25183) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24657) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24669) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17947), .QN(n24952) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24670) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24592) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17944), .QN(n24916) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n14401), .QN(n25105) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17943), .QN(n25269) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17942), .QN(n25279) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17941), .QN(n25097) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2140) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2136) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2137) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2133) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2126) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2134) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2123) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2124) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2120) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2121) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24735), .QN(n2127) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2118) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2142) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24595), .QN(n2143) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2139) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_5/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_5/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2117) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_5/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_5/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [5]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_5/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_5/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net366478), .QN(net740661) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_6/data_reg  ( .D(n23990), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17940) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_6/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_6/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_6/N3 ) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_6/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_6/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_6/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_6/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_6/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n17939) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24671) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17937), .QN(n25289) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17936), .QN(n25278) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17935), .QN(n24981) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17934), .QN(n25287) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24658) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24672) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17931), .QN(n24953) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24673) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24593) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17928), .QN(n24917) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n14127), .QN(n25106) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17927), .QN(n25270) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17926), .QN(n25280) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17925), .QN(n25285) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2104) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2100) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2101) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2097) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2090) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n23260), .QN(n2098) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2087) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2088) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2084) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2085) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24738), .QN(n2091) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2082) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2106) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24597), .QN(n2107) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2103) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_6/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_6/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2081) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_6/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_6/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [6]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_6/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_6/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n5729), .QN(n25346) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_7/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_7/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_7/N3 ), .QN(n17924) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_7/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_7/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_7/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_7/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_7/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n17923) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24659) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17921), .QN(n25258) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17920), .QN(n25048) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17919), .QN(n24982) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17918), .QN(n25184) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24661) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24660) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17915), .QN(n25042) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24662) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24589) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17912), .QN(n24918) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n14399), .QN(n24778) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17911), .QN(n24890) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17910), .QN(n24845) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17909), .QN(n25037) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2068) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2064) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2065) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2061) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24792), .QN(n2054) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2062) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2051) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2052) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2048) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2049) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24600), .QN(n2055) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2046) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2070) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24726), .QN(n2071) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2067) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_7/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_7/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2045) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_7/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_7/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [7]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_7/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_7/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net366191), .QN(net740717) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_8/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_8/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_8/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_8/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_8/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n17908) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24663) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17906), .QN(n25259) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17905), .QN(n25049) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17904), .QN(n24983) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17903), .QN(n25185) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24665) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24664) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17900), .QN(n25043) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24666) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24590) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17897), .QN(n24919) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n14400), .QN(n24779) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17896), .QN(n24891) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17895), .QN(n24846) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17894), .QN(n25038) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2032) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2028) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2029) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2025) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24790), .QN(n2018) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2026) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2015) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2016) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2012) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2013) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24598), .QN(n2019) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2010) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2034) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24724), .QN(n2035) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2031) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_8/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_8/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2009) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_8/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_8/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [8]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_8/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_8/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net741293), .QN(n17893) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_10/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_10/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_10/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_10/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_10/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17892) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17891), .QN(n25001) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17890), .QN(n25252) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17889), .QN(n25203) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17888), .QN(n24973) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17887), .QN(n25177) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24631) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24632) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17884), .QN(n25155) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17883), .QN(n25147) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17882), .QN(n25109) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17881), .QN(n24894) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17880), .QN(n25265) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17879), .QN(n25100) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17878), .QN(n25273) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17877), .QN(n24852) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3076) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3072) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3073) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3069) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3062) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3070) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3059) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3060) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24701), .QN(n3056) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3057) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3063) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24688), .QN(n3054) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24703), .QN(n3078) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24702), .QN(n3079) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3075) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_10/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3053) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_10/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_10/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [10]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_10/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_10/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24601), .QN(n4416) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_11/data_reg  ( .D(n11725), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17876) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_11/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_11/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_11/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_11/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_11/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17875) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17874), .QN(n25002) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17873), .QN(n25253) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17872), .QN(n25204) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17871), .QN(n24974) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17870), .QN(n25178) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24633) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24634) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17867), .QN(n25156) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17866), .QN(n25148) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17865), .QN(n25110) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17864), .QN(n24895) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17863), .QN(n25266) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17862), .QN(n25101) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17861), .QN(n25274) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17860), .QN(n24853) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3040) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3036) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3037) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3033) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3026) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3034) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3023) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3024) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24704), .QN(n3020) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3021) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3027) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24685), .QN(n3018) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24706), .QN(n3042) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24705), .QN(n3043) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3039) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_11/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3017) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_11/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_11/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [11]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_11/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_11/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24812), .QN(n17859) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_12/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_12/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_12/N3 ) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_12/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_12/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_12/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_12/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_12/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17858) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17857), .QN(n24822) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17856), .QN(n24829) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17855), .QN(n24828) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17854), .QN(n24821) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17853), .QN(n24827) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24620) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24621) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17850), .QN(n24826) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17849), .QN(n24825) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17848), .QN(n24824) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17847), .QN(n24820) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17846), .QN(n24842) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17845), .QN(n24823) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17844), .QN(n24831) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17843), .QN(n24819) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3004) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3000) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3001) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2997) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2990) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2998) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2987) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2988) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24682), .QN(n2984) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2985) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2991) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24681), .QN(n2982) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24684), .QN(n3006) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24683), .QN(n3007) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n3003) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_12/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_12/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2981) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_12/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_12/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [12]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_12/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_12/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24811), .QN(n4410) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_14/data_reg  ( .D(net767257), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17842) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_14/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_14/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_14/N3 ) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_14/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_14/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_14/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_14/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_14/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17841) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17840), .QN(n25004) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17839), .QN(n25255) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17838), .QN(n25206) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17837), .QN(n24976) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17836), .QN(n25180) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24637) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24638) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17833), .QN(n25158) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17832), .QN(n25150) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17831), .QN(n25112) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17830), .QN(n24897) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17829), .QN(n25267) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17828), .QN(n25103) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17827), .QN(n25275) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17826), .QN(n24855) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2932) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2928) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2929) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2925) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2918) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2926) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2915) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2916) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24709), .QN(n2912) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2913) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2919) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24690), .QN(n2910) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24711), .QN(n2934) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24710), .QN(n2935) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2931) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_14/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_14/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2909) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_14/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_14/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [14]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_14/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_14/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24814), .QN(n4404) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_15/data_reg  ( .D(n23986), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17825) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_15/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_15/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_15/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_15/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_15/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17824) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17823), .QN(n25005) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17822), .QN(n25256) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17821), .QN(n25207) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17820), .QN(n24977) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17819), .QN(n25181) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24639) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24640) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17816), .QN(n25159) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17815), .QN(n25151) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17814), .QN(n25113) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17813), .QN(n24898) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17812), .QN(n25268) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17811), .QN(n25104) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17810), .QN(n25276) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17809), .QN(n24856) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2896) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2892) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2893) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2889) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2882) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2890) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2879) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2880) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24712), .QN(n2876) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2877) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2883) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24689), .QN(n2874) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24714), .QN(n2898) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24713), .QN(n2899) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2895) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_15/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_15/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2873) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_15/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_15/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [15]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_15/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_15/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24810), .QN(n4401) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_13/data_reg  ( .D(n11847), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17808) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_13/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_13/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_13/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_13/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_13/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17807) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17806), .QN(n25003) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17805), .QN(n25254) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17804), .QN(n25205) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17803), .QN(n24975) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17802), .QN(n25179) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17801), .QN(n25174) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24635) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17799), .QN(n25157) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17798), .QN(n25149) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n14402), .QN(n25111) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17797), .QN(n24896) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17796), .QN(n25305) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17795), .QN(n25102) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17794), .QN(n24858) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17793), .QN(n24854) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24708), .QN(n2968) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24747), .QN(n2964) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2965) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24794), .QN(n2961) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2954) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2962) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2951) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n2952) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24707), .QN(n2948) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24636) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n998), .QN(n25078) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n997), .QN(n25046) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n996), .QN(n24875) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n995), .QN(n24859) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n994), .QN(n25081) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_13/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_13/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n993), .QN(n24847) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_13/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_13/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [13]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_13/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_13/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n991), .QN(n25347) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_16/data_reg  ( .D(
        \core_inst/IFID_NPC/DFF_16/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n17792) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_16/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_16/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_16/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_16/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_16/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17791) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17790), .QN(n25006) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24749), .QN(n983) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17789), .QN(n25208) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n981) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n980) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n979) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n978) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17788), .QN(n25160) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n23261), .QN(n976) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17787), .QN(n25114) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17786), .QN(n24899) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n973) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24748), .QN(n972) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24715), .QN(n971) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24729), .QN(n970) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n969), .QN(n25021) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n968), .QN(n25237) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n967), .QN(n25050) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n966), .QN(n25222) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n965), .QN(n25186) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n964), .QN(n24984) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n963), .QN(n24956) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24641) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n961), .QN(n24936) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n960), .QN(n25130) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n959), .QN(n24921) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n958), .QN(n25065) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n957), .QN(n24876) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n956), .QN(n24860) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n955), .QN(n25082) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_16/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_16/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n954), .QN(n25290) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_16/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_16/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n952), .QN(n25348) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_18/data_reg  ( .D(n23987), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17785) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_18/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_18/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_18/N3 ) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_18/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_18/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_18/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_18/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_18/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17784) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17783), .QN(n25008) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24740), .QN(n943) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17782), .QN(n25210) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n941) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n940) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n939) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n938) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17781), .QN(n25162) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n936) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17780), .QN(n25116) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17779), .QN(n24901) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n933) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24739), .QN(n932) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24691), .QN(n931) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24803), .QN(n930) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n929), .QN(n25023) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n928), .QN(n25239) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n927), .QN(n25052) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n926), .QN(n25224) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n925), .QN(n25188) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n924), .QN(n24986) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n923), .QN(n24958) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24622) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n921), .QN(n24938) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n920), .QN(n25132) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n919), .QN(n24923) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n918), .QN(n25067) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n917), .QN(n24878) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n916), .QN(n24862) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n915), .QN(n25084) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_18/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_18/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n914), .QN(n25292) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_18/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_18/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [18]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_18/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_18/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n912), .QN(n25283) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_19/data_reg  ( .D(net780182), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17778) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_19/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_19/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_19/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_19/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_19/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17777) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17776), .QN(n25009) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24753), .QN(n904) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17775), .QN(n25211) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n902) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n901) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n900) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n899) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17774), .QN(n25163) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n897) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17773), .QN(n25117) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17772), .QN(n24902) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n894) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24752), .QN(n893) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24717), .QN(n892) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24731), .QN(n891) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n890), .QN(n25024) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n889), .QN(n25240) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n888), .QN(n25053) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n887), .QN(n25225) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n886), .QN(n25189) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n885), .QN(n24987) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n884), .QN(n24959) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24643) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n882), .QN(n24939) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n881), .QN(n25133) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n880), .QN(n24924) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n879), .QN(n25068) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n878), .QN(n24879) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n877), .QN(n24863) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n876), .QN(n25085) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_19/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_19/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n875), .QN(n25293) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_19/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_19/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [19]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_19/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_19/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n873), .QN(n25308) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_20/data_reg  ( .D(n22840), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17771) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_20/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_20/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_20/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_20/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_20/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17770) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17769), .QN(net741056) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net741388), .QN(n865) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17768), .QN(net740836) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n863) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n862) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n861) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n860) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17767), .QN(net740888) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n858) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17766), .QN(net740938) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17765), .QN(net741172) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n855) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net741389), .QN(n854) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net741442), .QN(n853) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net741397), .QN(n852) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n851), .QN(net741039) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n850), .QN(net740803) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n849), .QN(net741008) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n848), .QN(net740820) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n847), .QN(net740860) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n846), .QN(net741080) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n845), .QN(net741110) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(net741520) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n843), .QN(net741132) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n842), .QN(net740920) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n841), .QN(net741149) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n840), .QN(net740991) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n839), .QN(net741198) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n838), .QN(net741216) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n837), .QN(net740972) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_20/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_20/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n836), .QN(net740741) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_20/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_20/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [20]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_20/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_20/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n834), .QN(n25309) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_22/data_reg  ( .D(n23983), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17764) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_22/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_22/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_22/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_22/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_22/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17763) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17762), .QN(net741054) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net741384), .QN(n825) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17761), .QN(net740834) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n823) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n822) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n821) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n820) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17760), .QN(net740886) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n818) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17759), .QN(net740936) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17758), .QN(net741170) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n815) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net741385), .QN(n814) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net741440), .QN(n813) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net741400), .QN(n812) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n811), .QN(net741037) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n810), .QN(net740801) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n809), .QN(net741006) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n808), .QN(net740818) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n807), .QN(net740858) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n806), .QN(net741078) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n805), .QN(net741108) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(net741518) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n803), .QN(net741130) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n802), .QN(net740918) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n801), .QN(net741147) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n800), .QN(net740989) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n799), .QN(net741196) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n798), .QN(net741214) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n797), .QN(net740970) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_22/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_22/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n796), .QN(net740739) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_22/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_22/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [22]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_22/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_22/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n794), .QN(net740721) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_23/data_reg  ( .D(n23991), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17757) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_23/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_23/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_23/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_23/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_23/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17756) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17755), .QN(n25011) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24755), .QN(n786) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17754), .QN(n25213) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n784) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n783) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n782) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n781) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17753), .QN(n25165) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n779) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17752), .QN(n25119) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17751), .QN(n24905) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n776) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24754), .QN(n775) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24718), .QN(n774) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24733), .QN(n773) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n772), .QN(n25026) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n771), .QN(n25242) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n770), .QN(n25055) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n769), .QN(n25227) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n768), .QN(n25191) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n767), .QN(n24989) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n766), .QN(n24961) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24644) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n764), .QN(n24941) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n763), .QN(n25135) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n762), .QN(n24926) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n761), .QN(n25070) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n760), .QN(n24881) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n759), .QN(n24865) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n758), .QN(n25087) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_23/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_23/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n757), .QN(n25295) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_23/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_23/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [23]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_23/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_23/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n755), .QN(n25311) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_21/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_21/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_21/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_21/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_21/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17750) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17749), .QN(n25010) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24742), .QN(n748) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17748), .QN(n25212) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n746) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n745) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n744) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n743) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17747), .QN(n25164) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n741) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17746), .QN(n25118) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17745), .QN(n24904) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n738) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24741), .QN(n737) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24692), .QN(n736) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24800), .QN(n735) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n734), .QN(n25025) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n733), .QN(n25241) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n732), .QN(n25054) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n731), .QN(n25226) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n730), .QN(n25190) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n729), .QN(n24988) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n728), .QN(n24960) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24624) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n726), .QN(n24940) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n725), .QN(n25134) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n724), .QN(n24925) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n723), .QN(n25069) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n722), .QN(n24880) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n721), .QN(n24864) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n720), .QN(n25086) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_21/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_21/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n719), .QN(n25294) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_21/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_21/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [21]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_21/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_21/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n717), .QN(n25307) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_17/data_reg  ( .D(n23985), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17744) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_17/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_17/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_17/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_17/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_17/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17742) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17741), .QN(n25007) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24751), .QN(n710) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17740), .QN(n25209) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n708) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n707) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n706) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n705) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17739), .QN(n25161) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n703) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17738), .QN(n25115) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17737), .QN(n24900) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n700) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24750), .QN(n699) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24716), .QN(n698) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24730), .QN(n697) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n696), .QN(n25022) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n695), .QN(n25238) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n694), .QN(n25051) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n693), .QN(n25223) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n692), .QN(n25187) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n691), .QN(n24985) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n690), .QN(n24957) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24642) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n688), .QN(n24937) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n687), .QN(n25131) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n686), .QN(n24922) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n685), .QN(n25066) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n684), .QN(n24877) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n683), .QN(n24861) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n682), .QN(n25083) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_17/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_17/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n681), .QN(n25291) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_17/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_17/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [17]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_17/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_17/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n679), .QN(n25312) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_24/data_reg  ( .D(n23984), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17736) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_24/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_24/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_24/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_24/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_24/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17735) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17734), .QN(n25012) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24757), .QN(n671) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17733), .QN(n25214) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n669) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n668) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n667) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n666) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17732), .QN(n25166) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n664) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17731), .QN(n25120) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17730), .QN(n24906) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n661) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24756), .QN(n660) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24719), .QN(n659) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24734), .QN(n658) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n657), .QN(n25027) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n656), .QN(n25243) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n655), .QN(n25056) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n654), .QN(n25228) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n653), .QN(n25192) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n652), .QN(n24990) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n651), .QN(n24962) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24645) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n649), .QN(n24942) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n648), .QN(n25136) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n647), .QN(n24927) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n646), .QN(n25071) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n645), .QN(n24882) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n644), .QN(n24866) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n643), .QN(n25088) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_24/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_24/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n642), .QN(n25296) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_24/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_24/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [24]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_24/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_24/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n640), .QN(net740655) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_26/data_reg  ( .D(n14058), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17729) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_26/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_26/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_26/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_26/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_26/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17728) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17727), .QN(n25014) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24744), .QN(n631) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17726), .QN(n25216) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n629) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n628) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n627) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n626) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17725), .QN(n25168) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n624) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17724), .QN(n25122) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17723), .QN(n24908) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n621) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24743), .QN(n620) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24693), .QN(n619) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24796), .QN(n618) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n617), .QN(n25029) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n616), .QN(n25245) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n615), .QN(n25058) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n614), .QN(n25230) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n613), .QN(n25194) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n612), .QN(n24992) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n611), .QN(n24964) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24625) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n609), .QN(n24944) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n608), .QN(n25138) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n607), .QN(n24929) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n606), .QN(n25073) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n605), .QN(n24884) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n604), .QN(n24868) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n603), .QN(n25090) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_26/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_26/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n602), .QN(n25298) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_26/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_26/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n600), .QN(n25350) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_27/data_reg  ( .D(n23980), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17722) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_27/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_27/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_27/N3 ) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_27/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_27/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_27/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_27/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_27/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17720) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17719), .QN(n25015) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24761), .QN(n592) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17718), .QN(n25217) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n590) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n589) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n588) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n587) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17717), .QN(n25169) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n585) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17716), .QN(n25123) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17715), .QN(n24909) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n582) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24760), .QN(n581) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24721), .QN(n580) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24797), .QN(n579) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n578), .QN(n25030) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n577), .QN(n25246) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n576), .QN(n25059) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n575), .QN(n25231) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n574), .QN(n25195) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n573), .QN(n24993) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n572), .QN(n24965) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24647) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n570), .QN(n24945) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n569), .QN(n25139) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n568), .QN(n24930) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n567), .QN(n25074) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n566), .QN(n24885) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n565), .QN(n24869) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n564), .QN(n25091) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_27/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_27/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n563), .QN(n25299) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_27/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_27/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [27]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_27/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_27/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n561), .QN(n25354) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_28/data_reg  ( .D(net812861), .CK(DLX_CLK), 
        .RN(DLX_RST), .QN(n22701) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_28/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_28/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_28/N3 ) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_28/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_28/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_28/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_28/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_28/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17713) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17712), .QN(n25016) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24763), .QN(n553) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17711), .QN(n25218) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n551) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n550) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n549) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n548) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17710), .QN(n25170) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n546) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17709), .QN(n25124) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17708), .QN(n24910) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n543) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24762), .QN(n542) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24722), .QN(n541) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24799), .QN(n540) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n539), .QN(n25031) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n538), .QN(n25247) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n537), .QN(n25060) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n536), .QN(n25232) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n535), .QN(n25196) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n534), .QN(n24994) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n533), .QN(n24966) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24648) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n531), .QN(n24946) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n530), .QN(n25140) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n529), .QN(n24931) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n528), .QN(n25075) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n527), .QN(n24886) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n526), .QN(n24870) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n525), .QN(n25092) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_28/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_28/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n524), .QN(n25300) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_28/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_28/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n522) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_30/data_reg  ( .D(n23989), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17707) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_30/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_30/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_30/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_30/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_30/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17706) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17705), .QN(n25018) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24765), .QN(n513) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17704), .QN(n25220) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n511) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n510) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n509) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n508) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17703), .QN(n25172) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n506) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17702), .QN(n25126) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17701), .QN(n24913) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n503) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24764), .QN(n502) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24723), .QN(n501) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24795), .QN(n500) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n499), .QN(n25033) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n498), .QN(n25249) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n497), .QN(n25062) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n496), .QN(n25234) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n495), .QN(n25198) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n494), .QN(n24996) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n493), .QN(n24968) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24653) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n491), .QN(n24948) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n490), .QN(n25142) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n489), .QN(n24933) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n488), .QN(n25077) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n487), .QN(n24888) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n486), .QN(n24872) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n485), .QN(n25094) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_30/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_30/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n484), .QN(n25302) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_30/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_30/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [30]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_30/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_30/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n482), .QN(n25349) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_31/data_reg  ( .D(n23992), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17700) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_31/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_31/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_31/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_31/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_31/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17699) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n475) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n474) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n473) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n472) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24766), .QN(n471) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24767), .QN(n470) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24768), .QN(n469) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n468) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17698), .QN(n25127) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17697), .QN(n24914) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n465) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24769), .QN(n464) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n463) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24798), .QN(n462) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n461), .QN(n25034) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24656) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n459), .QN(n25063) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n458), .QN(n25235) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n457), .QN(n25199) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n456), .QN(n24997) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n455), .QN(n24969) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n454), .QN(n24954) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n453), .QN(n24949) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n452), .QN(n25143) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n451), .QN(n24934) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24654) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24655) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n448), .QN(n24873) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n447), .QN(n25095) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_31/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_31/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n446), .QN(n24848) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_29/data_reg  ( .D(n23988), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17696) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_29/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_29/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_29/N3 ) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_29/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_29/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_29/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_29/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_29/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17695) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17694), .QN(n25017) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24746), .QN(n439) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17693), .QN(n25219) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n437) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n436) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n435) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n434) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17692), .QN(n25171) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n432) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17691), .QN(n25125) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17690), .QN(n24911) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n429) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24745), .QN(n428) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24694), .QN(n427) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24802), .QN(n426) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n425), .QN(n25032) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n424), .QN(n25248) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n423), .QN(n25061) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n422), .QN(n25233) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n421), .QN(n25197) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n420), .QN(n24995) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n419), .QN(n24967) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24626) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n417), .QN(n24947) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n416), .QN(n25141) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n415), .QN(n24932) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n414), .QN(n25076) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n413), .QN(n24887) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n412), .QN(n24871) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n411), .QN(n25093) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_29/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_29/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n410), .QN(n25301) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_29/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_29/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [29]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_29/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_29/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24817), .QN(n4356) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_25/data_reg  ( .D(n23982), .CK(DLX_CLK), 
        .RN(DLX_RST), .QN(n17689) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_25/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_25/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_25/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_25/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_25/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17688) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17687), .QN(n25013) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24759), .QN(n401) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17686), .QN(n25215) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n399) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n398) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n397) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n396) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17685), .QN(n25167) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n394) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17684), .QN(n25121) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17683), .QN(n24907) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n391) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24758), .QN(n390) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24720), .QN(n389) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24732), .QN(n388) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n387), .QN(n25028) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n386), .QN(n25244) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n385), .QN(n25057) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n384), .QN(n25229) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n383), .QN(n25193) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n382), .QN(n24991) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n381), .QN(n24963) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24646) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n379), .QN(n24943) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n378), .QN(n25137) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n377), .QN(n24928) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n376), .QN(n25072) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n375), .QN(n24883) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n374), .QN(n24867) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n373), .QN(n25089) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_25/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_25/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n372), .QN(n25297) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_25/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_25/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [25]) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_25/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_25/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n24816), .QN(n4368) );
  DFFR_X1 \core_inst/EXMEM_NPC/DFF_9/data_reg  ( .D(
        \core_inst/EXMEM_NPC/DFF_9/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_NPC/DFF_9/N3 ) );
  DFFR_X1 \core_inst/MEMWB_NPC/DFF_9/data_reg  ( .D(
        \core_inst/MEMWB_NPC/DFF_9/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n17682) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_8/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17681), .QN(n25020) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_7/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n363) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_31/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17680), .QN(n25221) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_29/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n361) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_28/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n360) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_27/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24770), .QN(n359) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_26/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24771), .QN(n358) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_23/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17679), .QN(n25173) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_22/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n356) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_18/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17678), .QN(n25129) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_17/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n17677), .QN(n24920) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_16/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n353) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_15/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24772), .QN(n352) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_12/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n351) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_11/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n24801), .QN(n350) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_9/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n349), .QN(n25035) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_6/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n348), .QN(n25079) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_5/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n347), .QN(n25064) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_4/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n346), .QN(n25236) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_30/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n345), .QN(n25200) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_3/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n344), .QN(n24998) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_25/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n343), .QN(n24970) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_24/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n342), .QN(n24955) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_21/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n341), .QN(n24950) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_20/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n340), .QN(n25144) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_2/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n339), .QN(n24935) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_19/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n24667) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_14/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n337), .QN(n25303) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_13/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n336), .QN(n24874) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_10/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n335), .QN(n25096) );
  DFFR_X1 \core_inst/ID/REGISTER_FILE/REG_1/DFF_9/data_reg  ( .D(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_9/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n334), .QN(n24849) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_9/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_9/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n5761), .QN(n25310) );
  TBUF_X2 \core_inst/s_DRAM_DLX_OUT_tri[7]  ( .A(DRAM_INTERFACE[7]), .EN(n298), 
        .Z(\core_inst/MEM/MUX_LOAD/MUX_BIT_7/s_top ) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_29/data_reg  ( .D(
        \core_inst/IDEX_IR/DFF_29/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n14130), 
        .QN(net718078) );
  DFFR_X1 \core_inst/EXMEM_IR/DFF_27/data_reg  ( .D(
        \core_inst/EXMEM_IR/DFF_27/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n11743), .QN(n24574) );
  DFFR_X1 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_9/data_reg  ( .D(n16391), 
        .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [9]), .QN(n6460) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_27/data_reg  ( .D(
        \core_inst/IDEX_IR/DFF_27/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n15079), 
        .QN(net741262) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_4/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_4/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n25352) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_14/data_reg  ( .D(n22831), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n22736), .QN(n25323) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_8/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_8/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n5609) );
  DFFR_X1 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_10/data_reg  ( .D(
        \core_inst/IF_stage/PROGRAM_COUNTER/DFF_10/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [10]) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_2/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_2/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net717454), .QN(n5601) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_0/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_0/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_0/N3 ) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_31/data_reg  ( .D(n22803), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17670), .QN(n22739) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_29/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_29/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n25333), .QN(n5596) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_24/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_24/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n5595) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_22/data_reg  ( .D(n22719), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n24526), .QN(n25320) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_10/data_reg  ( .D(n22705), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n17665) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_3/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n5589) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_13/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_13/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_13/N3 ) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_10/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_10/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_10/N3 ) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_6/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_6/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17663) );
  DFFR_X1 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_7/data_reg  ( .D(net522736), 
        .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [7]), .QN(n5576) );
  DFFR_X1 \core_inst/IFID_IR/DFF_14/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_14/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(n6562)
         );
  DFFR_X1 \core_inst/MEMWB_IR/DFF_27/data_reg  ( .D(n24316), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(s_MEMWB_IR[27]), .QN(net718139) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_13/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_13/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n22946), .QN(n5186) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_10/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_10/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n25357) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_29/data_reg  ( .D(n22730), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n25351) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_26/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_26/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [26]) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_16/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_16/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [16]) );
  DFFR_X1 \core_inst/EXMEM_DATAIN/DFF_28/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_28/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/ps_EXMEM_DATA_IN [28]) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_12/data_reg  ( .D(net712313), .CK(DLX_CLK), .RN(DLX_RST), .QN(net89402) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_13/data_reg  ( .D(n26742), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n1660) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_2/data_reg  ( .D(n15062), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n6475) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_0/data_reg  ( .D(n22824), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n22732) );
  DFFR_X1 \core_inst/MEMWB_IR/DFF_26/data_reg  ( .D(n14429), .CK(DLX_CLK), 
        .RN(DLX_RST), .QN(net749529) );
  DFFR_X1 \core_inst/MEMWB_DATAOUT/DFF_3/data_reg  ( .D(
        \core_inst/MEMWB_DATAOUT/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n5307), .QN(net741572) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_30/data_reg  ( .D(
        \core_inst/IDEX_IR/DFF_30/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n14389), 
        .QN(net718077) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_25/data_reg  ( .D(n26781), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net366411), .QN(n25592) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_14/data_reg  ( .D(n26743), .CK(DLX_CLK), 
        .RN(DLX_RST), .QN(n6330) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_26/data_reg  ( .D(
        \core_inst/IDEX_IR/DFF_26/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        net741576) );
  DFFR_X1 \cu_inst/WB/DFF_3/data_reg  ( .D(\cu_inst/WB/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(s_ID_rf_write_en) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_9/data_reg  ( .D(n22938), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n6555) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_21/data_reg  ( .D(n22841), .CK(DLX_CLK), 
        .RN(DLX_RST), .QN(n753) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_19/data_reg  ( .D(n22740), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net718081), .QN(n1668) );
  DFFS_X1 \core_inst/EXMEM_IR/DFF_28/data_reg  ( .D(n13343), .CK(DLX_CLK), 
        .SN(DLX_RST), .Q(\cu_inst/FW_UNIT/ITD_EXMEM/N17 ), .QN(n25581) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_7/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_7/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n5618) );
  DFFS_X2 \cu_inst/MEM/DFF_7/data_reg  ( .D(n1600), .CK(DLX_CLK), .SN(DLX_RST), 
        .Q(n298), .QN(\core_inst/N65 ) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_20/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_20/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n5187) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_9/data_reg  ( .D(n22731), .CK(DLX_CLK), 
        .RN(DLX_RST), .QN(n25360) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_23/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_23/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n25363) );
  DFFR_X1 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_11/data_reg  ( .D(
        \core_inst/IF_stage/PROGRAM_COUNTER/DFF_11/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [11]), .QN(n5577) );
  DFFR_X1 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_26/data_reg  ( .D(n26783), 
        .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [26]) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_21/data_reg  ( .D(n22825), .CK(DLX_CLK), 
        .RN(DLX_RST), .QN(n716) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_22/data_reg  ( .D(n22852), .CK(DLX_CLK), 
        .RN(DLX_RST), .QN(n793) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_0/data_reg  ( .D(n22706), .CK(DLX_CLK), 
        .RN(DLX_RST), .QN(n1537) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_27/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_27/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n562) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_19/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_19/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        net740632) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_24/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_24/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n25340) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_10/data_reg  ( .D(n22707), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n22823), .QN(n1187) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_27/data_reg  ( .D(n22806), .CK(DLX_CLK), 
        .RN(DLX_RST), .Q(n14769) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_8/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_8/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n25322) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_13/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_13/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n25355) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_23/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_23/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n22802), .QN(n756) );
  DFFS_X1 \core_inst/MEMWB_IR/DFF_18/data_reg  ( .D(n1649), .CK(DLX_CLK), .SN(
        DLX_RST), .Q(n25591), .QN(s_MEMWB_IR[18]) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_5/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_5/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n22942), .QN(n25321) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_16/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_16/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n953) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_10/data_reg  ( .D(n22843), .CK(DLX_CLK), 
        .RN(DLX_RST), .QN(n1222) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_7/data_reg  ( .D(n22815), .CK(DLX_CLK), .RN(
        DLX_RST), .QN(n1301) );
  DFFR_X1 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_19/data_reg  ( .D(n16388), 
        .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [19]), .QN(n6512) );
  NAND3_X1 U15863 ( .A1(s_IFID_IR[17]), .A2(s_IFID_IR[19]), .A3(net741547), 
        .ZN(n19261) );
  NAND3_X1 U15864 ( .A1(s_IFID_IR[18]), .A2(s_IFID_IR[17]), .A3(net741696), 
        .ZN(n19249) );
  NAND3_X1 U15884 ( .A1(s_IFID_IR[24]), .A2(s_IFID_IR[22]), .A3(n24582), .ZN(
        n20080) );
  NAND3_X1 U15885 ( .A1(s_IFID_IR[23]), .A2(s_IFID_IR[22]), .A3(n24586), .ZN(
        n20070) );
  NAND3_X1 U15886 ( .A1(s_IFID_IR[23]), .A2(s_IFID_IR[24]), .A3(n24618), .ZN(
        n20065) );
  NAND3_X1 U15887 ( .A1(n24586), .A2(n24582), .A3(n24618), .ZN(n20081) );
  NAND3_X1 U15891 ( .A1(n20118), .A2(n18153), .A3(n18179), .ZN(n18143) );
  DFFRS_X1 \core_inst/IDEX_RF_ADDR_DEST/DFF_3/data_reg  ( .D(
        \core_inst/IDEX_RF_ADDR_DEST/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), 
        .SN(1'b1), .Q(n17654) );
  DFFRS_X1 \core_inst/IDEX_RF_ADDR_DEST/DFF_4/data_reg  ( .D(
        \core_inst/IDEX_RF_ADDR_DEST/DFF_4/N3 ), .CK(DLX_CLK), .RN(DLX_RST), 
        .SN(1'b1), .Q(n17656) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_17/data_reg  ( .D(n22810), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net718082), .QN(n1666) );
  DFFR_X1 \core_inst/IDEX_IR/DFF_16/data_reg  ( .D(n22828), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(net718086), .QN(n1665) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[0]  ( .A(n297), .EN(n298), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_0/s_top ) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[0]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_0/s_top ), .EN(\core_inst/N65 ), .Z(
        DRAM_INTERFACE[0]) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[0]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [0]), .EN(\core_inst/N65 ), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_0/s_top ) );
  DFFR_X1 \cu_inst/EX/DFF_10/data_reg  ( .D(\cu_inst/EX/DFF_10/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(s_EX_BOT_MUX), .QN(net740706) );
  DFFR_X2 \cu_inst/EX/DFF_17/data_reg  ( .D(\cu_inst/EX/DFF_17/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(net366451), .QN(net741458) );
  DFFRS_X1 \core_inst/IDEX_RF_ADDR_DEST/DFF_2/data_reg  ( .D(
        \core_inst/IDEX_RF_ADDR_DEST/DFF_2/N3 ), .CK(DLX_CLK), .RN(DLX_RST), 
        .SN(1'b1), .Q(n17657) );
  DFFRS_X1 \core_inst/IDEX_RF_ADDR_DEST/DFF_0/data_reg  ( .D(
        \core_inst/IDEX_RF_ADDR_DEST/DFF_0/N3 ), .CK(DLX_CLK), .RN(DLX_RST), 
        .SN(1'b1), .QN(n22674) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_8/data_reg  ( .D(n22947), .CK(DLX_CLK), .RN(
        DLX_RST), .Q(n13824) );
  DFFR_X1 \core_inst/IFID_NPC/DFF_12/data_reg  ( .D(
        \core_inst/IFID_NPC/DFF_12/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n13778) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[22]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[22] ), .EN(n25684), .Z(DRAM_INTERFACE[22])
         );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[23]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[23] ), .EN(n25684), .Z(DRAM_INTERFACE[23])
         );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[21]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[21] ), .EN(n25684), .Z(DRAM_INTERFACE[21])
         );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[20]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[20] ), .EN(n25684), .Z(DRAM_INTERFACE[20])
         );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[19]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[19] ), .EN(n25684), .Z(DRAM_INTERFACE[19])
         );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[18]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[18] ), .EN(n25684), .Z(DRAM_INTERFACE[18])
         );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[17]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[17] ), .EN(n25684), .Z(DRAM_INTERFACE[17])
         );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[16]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[16] ), .EN(n25684), .Z(DRAM_INTERFACE[16])
         );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[15]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_15/s_top ), .EN(n25684), .Z(
        DRAM_INTERFACE[15]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[14]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_14/s_top ), .EN(n25684), .Z(
        DRAM_INTERFACE[14]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[13]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_13/s_top ), .EN(n25684), .Z(
        DRAM_INTERFACE[13]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[12]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_12/s_top ), .EN(n25684), .Z(
        DRAM_INTERFACE[12]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[11]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_11/s_top ), .EN(n25684), .Z(
        DRAM_INTERFACE[11]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[10]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_10/s_top ), .EN(n25684), .Z(
        DRAM_INTERFACE[10]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[9]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_9/s_top ), .EN(n25684), .Z(
        DRAM_INTERFACE[9]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[8]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_8/s_top ), .EN(n25684), .Z(
        DRAM_INTERFACE[8]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[6]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_6/s_top ), .EN(n25684), .Z(
        DRAM_INTERFACE[6]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[5]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_5/s_top ), .EN(n25684), .Z(
        DRAM_INTERFACE[5]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[4]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_4/s_top ), .EN(n25684), .Z(
        DRAM_INTERFACE[4]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[3]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_3/s_top ), .EN(n25684), .Z(
        DRAM_INTERFACE[3]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[2]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_2/s_top ), .EN(n25684), .Z(
        DRAM_INTERFACE[2]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[1]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_1/s_top ), .EN(n25684), .Z(
        DRAM_INTERFACE[1]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[31]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[31] ), .EN(\core_inst/N65 ), .Z(
        DRAM_INTERFACE[31]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[30]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[30] ), .EN(\core_inst/N65 ), .Z(
        DRAM_INTERFACE[30]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[29]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[29] ), .EN(\core_inst/N65 ), .Z(
        DRAM_INTERFACE[29]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[28]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[28] ), .EN(\core_inst/N65 ), .Z(
        DRAM_INTERFACE[28]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[27]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[27] ), .EN(\core_inst/N65 ), .Z(
        DRAM_INTERFACE[27]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[26]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[26] ), .EN(\core_inst/N65 ), .Z(
        DRAM_INTERFACE[26]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[25]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[25] ), .EN(\core_inst/N65 ), .Z(
        DRAM_INTERFACE[25]) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[24]  ( .A(
        \core_inst/s_DRAM_DLX_OUT[24] ), .EN(\core_inst/N65 ), .Z(
        DRAM_INTERFACE[24]) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[6]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [6]), .EN(n25684), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_6/s_top ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[5]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [5]), .EN(n25684), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_5/s_top ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[4]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [4]), .EN(n25684), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_4/s_top ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[3]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [3]), .EN(n25684), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_3/s_top ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[2]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [2]), .EN(n25684), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_2/s_top ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[1]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [1]), .EN(n25684), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_1/s_top ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[6]  ( .A(DRAM_INTERFACE[6]), .EN(n298), 
        .Z(\core_inst/MEM/MUX_LOAD/MUX_BIT_6/s_top ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[5]  ( .A(DRAM_INTERFACE[5]), .EN(n298), 
        .Z(\core_inst/MEM/MUX_LOAD/MUX_BIT_5/s_top ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[4]  ( .A(DRAM_INTERFACE[4]), .EN(n298), 
        .Z(\core_inst/MEM/MUX_LOAD/MUX_BIT_4/s_top ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[3]  ( .A(DRAM_INTERFACE[3]), .EN(n298), 
        .Z(\core_inst/MEM/MUX_LOAD/MUX_BIT_3/s_top ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[2]  ( .A(DRAM_INTERFACE[2]), .EN(n298), 
        .Z(\core_inst/MEM/MUX_LOAD/MUX_BIT_2/s_top ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[1]  ( .A(DRAM_INTERFACE[1]), .EN(n298), 
        .Z(\core_inst/MEM/MUX_LOAD/MUX_BIT_1/s_top ) );
  DFFR_X1 \core_inst/IDEX_IMM_IN/DFF_7/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_7/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n24786) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[13]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [13]), .EN(n25684), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_13/s_top ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[11]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [11]), .EN(n25684), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_11/s_top ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[10]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [10]), .EN(n25684), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_10/s_top ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[13]  ( .A(DRAM_INTERFACE[13]), .EN(
        n298), .Z(\core_inst/MEM/MUX_LOAD/MUX_BIT_13/s_top ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[11]  ( .A(DRAM_INTERFACE[11]), .EN(
        n298), .Z(\core_inst/MEM/MUX_LOAD/MUX_BIT_11/s_top ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[10]  ( .A(DRAM_INTERFACE[10]), .EN(
        n298), .Z(\core_inst/MEM/MUX_LOAD/MUX_BIT_10/s_top ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[15]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [15]), .EN(n25684), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_15/s_top ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[15]  ( .A(DRAM_INTERFACE[15]), .EN(
        n298), .Z(\core_inst/MEM/MUX_LOAD/MUX_BIT_15/s_top ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[14]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [14]), .EN(n25684), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_14/s_top ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[12]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [12]), .EN(n25684), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_12/s_top ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[9]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [9]), .EN(n25684), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_9/s_top ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[8]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [8]), .EN(n25684), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_8/s_top ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[14]  ( .A(DRAM_INTERFACE[14]), .EN(
        n298), .Z(\core_inst/MEM/MUX_LOAD/MUX_BIT_14/s_top ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[12]  ( .A(DRAM_INTERFACE[12]), .EN(
        n298), .Z(\core_inst/MEM/MUX_LOAD/MUX_BIT_12/s_top ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[9]  ( .A(DRAM_INTERFACE[9]), .EN(n298), 
        .Z(\core_inst/MEM/MUX_LOAD/MUX_BIT_9/s_top ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[8]  ( .A(DRAM_INTERFACE[8]), .EN(n298), 
        .Z(\core_inst/MEM/MUX_LOAD/MUX_BIT_8/s_top ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[31]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [31]), .EN(n25684), .Z(
        \core_inst/s_DRAM_DLX_OUT[31] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[28]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [28]), .EN(\core_inst/N65 ), .Z(
        \core_inst/s_DRAM_DLX_OUT[28] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[17]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [17]), .EN(\core_inst/N65 ), .Z(
        \core_inst/s_DRAM_DLX_OUT[17] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[31]  ( .A(DRAM_INTERFACE[31]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[31] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[28]  ( .A(DRAM_INTERFACE[28]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[28] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[17]  ( .A(DRAM_INTERFACE[17]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[17] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[30]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [30]), .EN(\core_inst/N65 ), .Z(
        \core_inst/s_DRAM_DLX_OUT[30] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[29]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [29]), .EN(\core_inst/N65 ), .Z(
        \core_inst/s_DRAM_DLX_OUT[29] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[27]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [27]), .EN(\core_inst/N65 ), .Z(
        \core_inst/s_DRAM_DLX_OUT[27] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[26]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [26]), .EN(\core_inst/N65 ), .Z(
        \core_inst/s_DRAM_DLX_OUT[26] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[25]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [25]), .EN(\core_inst/N65 ), .Z(
        \core_inst/s_DRAM_DLX_OUT[25] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[24]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [24]), .EN(\core_inst/N65 ), .Z(
        \core_inst/s_DRAM_DLX_OUT[24] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[23]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [23]), .EN(\core_inst/N65 ), .Z(
        \core_inst/s_DRAM_DLX_OUT[23] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[22]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [22]), .EN(\core_inst/N65 ), .Z(
        \core_inst/s_DRAM_DLX_OUT[22] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[21]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [21]), .EN(\core_inst/N65 ), .Z(
        \core_inst/s_DRAM_DLX_OUT[21] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[20]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [20]), .EN(\core_inst/N65 ), .Z(
        \core_inst/s_DRAM_DLX_OUT[20] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[19]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [19]), .EN(\core_inst/N65 ), .Z(
        \core_inst/s_DRAM_DLX_OUT[19] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[18]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [18]), .EN(\core_inst/N65 ), .Z(
        \core_inst/s_DRAM_DLX_OUT[18] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[16]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [16]), .EN(\core_inst/N65 ), .Z(
        \core_inst/s_DRAM_DLX_OUT[16] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[30]  ( .A(DRAM_INTERFACE[30]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[30] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[29]  ( .A(DRAM_INTERFACE[29]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[29] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[27]  ( .A(DRAM_INTERFACE[27]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[27] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[26]  ( .A(DRAM_INTERFACE[26]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[26] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[25]  ( .A(DRAM_INTERFACE[25]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[25] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[24]  ( .A(DRAM_INTERFACE[24]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[24] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[23]  ( .A(DRAM_INTERFACE[23]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[23] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[22]  ( .A(DRAM_INTERFACE[22]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[22] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[21]  ( .A(DRAM_INTERFACE[21]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[21] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[20]  ( .A(DRAM_INTERFACE[20]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[20] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[19]  ( .A(DRAM_INTERFACE[19]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[19] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[18]  ( .A(DRAM_INTERFACE[18]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[18] ) );
  TBUF_X1 \core_inst/s_DRAM_DLX_OUT_tri[16]  ( .A(DRAM_INTERFACE[16]), .EN(
        n298), .Z(\core_inst/s_DRAM_DLX_OUT[16] ) );
  TBUF_X1 \core_inst/MEM/MEM_INTERFACE_tri[7]  ( .A(
        \core_inst/ps_EXMEM_DATA_IN [7]), .EN(\core_inst/N65 ), .Z(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_7/s_top ) );
  DFFR_X1 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_13/data_reg  ( .D(n26784), 
        .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [13]), .QN(n11848) );
  TBUF_X1 \core_inst/CORE_DRAM_INTERFACE_tri[7]  ( .A(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_7/s_top ), .EN(n25684), .Z(
        DRAM_INTERFACE[7]) );
  NOR3_X1 U12213 ( .A1(s_IFID_IR[29]), .A2(n14191), .A3(n24581), .ZN(n20117)
         );
  NOR4_X1 U12187 ( .A1(s_IFID_IR[29]), .A2(s_IFID_IR[27]), .A3(n14191), .A4(
        n24611), .ZN(n20049) );
  NAND2_X1 U12186 ( .A1(n19282), .A2(n24581), .ZN(n18171) );
  NAND2_X1 U12199 ( .A1(s_IFID_IR[26]), .A2(net741565), .ZN(n18138) );
  NOR4_X1 U12196 ( .A1(n24581), .A2(n24583), .A3(n24612), .A4(s_IFID_IR[28]), 
        .ZN(n18175) );
  NAND4_X1 U12190 ( .A1(n24581), .A2(n24583), .A3(net741565), .A4(n14191), 
        .ZN(n18132) );
  NAND4_X1 U12097 ( .A1(s_IFID_IR[28]), .A2(s_IFID_IR[29]), .A3(n24581), .A4(
        n24612), .ZN(n18153) );
  NAND2_X1 U12094 ( .A1(s_IFID_IR[28]), .A2(n20117), .ZN(n18172) );
  NOR2_X1 U12093 ( .A1(s_IFID_IR[26]), .A2(net741565), .ZN(n18166) );
  AOI22_X1 U12091 ( .A1(n18166), .A2(n20049), .B1(n24813), .B2(net741565), 
        .ZN(n18154) );
  OAI211_X1 U12090 ( .C1(net741565), .C2(n18172), .A(n18154), .B(n18171), .ZN(
        n18196) );
  NOR3_X1 U12079 ( .A1(n14128), .A2(n18188), .A3(n20111), .ZN(n18182) );
  NOR2_X1 U12077 ( .A1(n18182), .A2(n18181), .ZN(n18140) );
  NAND4_X1 U12075 ( .A1(n14195), .A2(n18059), .A3(n24785), .A4(n24585), .ZN(
        n18170) );
  NOR3_X1 U12073 ( .A1(n14210), .A2(n14190), .A3(n20111), .ZN(n18161) );
  AOI21_X1 U12069 ( .B1(n24616), .B2(n18059), .A(n20107), .ZN(n18187) );
  NOR3_X1 U12068 ( .A1(n24585), .A2(n24677), .A3(n18187), .ZN(n18145) );
  NOR3_X1 U12045 ( .A1(s_IFID_IR[24]), .A2(s_IFID_IR[23]), .A3(n24618), .ZN(
        n20084) );
  NAND2_X1 U12033 ( .A1(n20084), .A2(n20078), .ZN(n19326) );
  NOR3_X1 U12047 ( .A1(s_IFID_IR[24]), .A2(s_IFID_IR[22]), .A3(n24582), .ZN(
        n20077) );
  NAND2_X1 U12039 ( .A1(n20062), .A2(n20077), .ZN(n19383) );
  NAND2_X1 U12041 ( .A1(n20084), .A2(n20062), .ZN(n19395) );
  NAND2_X1 U12025 ( .A1(n20077), .A2(n20078), .ZN(n19366) );
  NAND2_X1 U12022 ( .A1(n20076), .A2(n20084), .ZN(n19367) );
  NOR3_X1 U12009 ( .A1(n24586), .A2(n24582), .A3(n24618), .ZN(n20071) );
  NOR3_X1 U11992 ( .A1(s_IFID_IR[23]), .A2(s_IFID_IR[22]), .A3(n24586), .ZN(
        n20063) );
  NAND2_X1 U11988 ( .A1(n20063), .A2(n20078), .ZN(n19370) );
  NAND2_X1 U11987 ( .A1(n20076), .A2(n20077), .ZN(n19365) );
  NAND2_X1 U11984 ( .A1(n20071), .A2(n20061), .ZN(n19390) );
  NAND2_X1 U11974 ( .A1(n20061), .A2(n20064), .ZN(n19389) );
  NAND2_X1 U11972 ( .A1(n20062), .A2(n20063), .ZN(n19378) );
  NAND2_X1 U11971 ( .A1(n20060), .A2(n20061), .ZN(n19388) );
  NAND2_X1 U11979 ( .A1(n20061), .A2(n20063), .ZN(n19384) );
  AOI22_X1 U11962 ( .A1(s_IFID_IR[21]), .A2(n19294), .B1(n26780), .B2(
        net741353), .ZN(n20041) );
  NOR3_X1 U11129 ( .A1(s_IFID_IR[17]), .A2(s_IFID_IR[19]), .A3(net741547), 
        .ZN(n19256) );
  NAND2_X1 U11124 ( .A1(n19265), .A2(n19240), .ZN(n18400) );
  NAND2_X1 U11128 ( .A1(n19239), .A2(n19256), .ZN(n18390) );
  NAND2_X1 U11116 ( .A1(n19265), .A2(n19257), .ZN(n18318) );
  NOR3_X1 U11078 ( .A1(s_IFID_IR[17]), .A2(s_IFID_IR[18]), .A3(net741696), 
        .ZN(n19241) );
  NAND2_X1 U11066 ( .A1(n19239), .A2(n19241), .ZN(n18388) );
  NAND2_X1 U11061 ( .A1(n19239), .A2(n19242), .ZN(n18394) );
  NAND2_X1 U11059 ( .A1(n19240), .A2(n19241), .ZN(n18382) );
  NAND2_X1 U11058 ( .A1(n19238), .A2(n19239), .ZN(n18393) );
  NAND2_X1 U11080 ( .A1(n19238), .A2(n19257), .ZN(n18367) );
  NAND2_X1 U11074 ( .A1(n19241), .A2(n19257), .ZN(n18369) );
  NAND2_X1 U11073 ( .A1(n19255), .A2(n19256), .ZN(n18361) );
  NAND2_X1 U11109 ( .A1(n19256), .A2(n19257), .ZN(n18362) );
  NAND2_X1 U11107 ( .A1(n19255), .A2(n19265), .ZN(n18363) );
  NAND2_X1 U11070 ( .A1(n19250), .A2(n19239), .ZN(n18395) );
  OAI22_X1 U10696 ( .A1(n784), .A2(n18315), .B1(n783), .B2(n18316), .ZN(n18794) );
  AOI22_X1 U10695 ( .A1(net767173), .A2(n767), .B1(n18321), .B2(n769), .ZN(
        n18796) );
  NAND2_X1 U10694 ( .A1(n18529), .A2(n761), .ZN(n18797) );
  OAI211_X1 U10693 ( .C1(n776), .C2(net518461), .A(n18796), .B(n18797), .ZN(
        n18795) );
  AOI211_X1 U10692 ( .C1(n18312), .C2(n770), .A(n18794), .B(n18795), .ZN(
        n18787) );
  AOI22_X1 U10698 ( .A1(n18307), .A2(n17755), .B1(net716405), .B2(n17754), 
        .ZN(n18801) );
  AOI22_X1 U10699 ( .A1(net767239), .A2(n24718), .B1(n18306), .B2(n771), .ZN(
        n18800) );
  AOI22_X1 U10700 ( .A1(n18310), .A2(n772), .B1(n18311), .B2(n758), .ZN(n18799) );
  AOI22_X1 U10691 ( .A1(net716461), .A2(n762), .B1(n18347), .B2(n768), .ZN(
        n18788) );
  NOR2_X1 U10689 ( .A1(n782), .A2(net767232), .ZN(n18791) );
  OAI22_X1 U10688 ( .A1(n781), .A2(net767237), .B1(net716477), .B2(n24644), 
        .ZN(n18792) );
  AOI211_X1 U10687 ( .C1(n757), .C2(n18343), .A(n18791), .B(n18792), .ZN(
        n18790) );
  AOI22_X1 U10690 ( .A1(n18338), .A2(n766), .B1(n18339), .B2(n763), .ZN(n18789) );
  AOI22_X1 U10704 ( .A1(n18330), .A2(n764), .B1(n18331), .B2(n17752), .ZN(
        n18804) );
  AOI22_X1 U10702 ( .A1(net767167), .A2(n759), .B1(n18326), .B2(n24754), .ZN(
        n18806) );
  AOI22_X1 U10701 ( .A1(n18300), .A2(n760), .B1(net767235), .B2(n24755), .ZN(
        n18798) );
  AOI22_X1 U10703 ( .A1(n18328), .A2(n17751), .B1(net767214), .B2(n17753), 
        .ZN(n18805) );
  OAI22_X1 U10608 ( .A1(n590), .A2(n18315), .B1(n589), .B2(n18316), .ZN(n18686) );
  AOI22_X1 U10607 ( .A1(net767173), .A2(n573), .B1(n18321), .B2(n575), .ZN(
        n18688) );
  NAND2_X1 U10606 ( .A1(n18529), .A2(n567), .ZN(n18689) );
  OAI211_X1 U10605 ( .C1(n582), .C2(net518461), .A(n18688), .B(n18689), .ZN(
        n18687) );
  AOI211_X1 U10604 ( .C1(n18312), .C2(n576), .A(n18686), .B(n18687), .ZN(
        n18679) );
  AOI22_X1 U10610 ( .A1(n18307), .A2(n17719), .B1(net716405), .B2(n17718), 
        .ZN(n18693) );
  AOI22_X1 U10611 ( .A1(net767239), .A2(n24721), .B1(n18306), .B2(n577), .ZN(
        n18692) );
  AOI22_X1 U10612 ( .A1(n18310), .A2(n578), .B1(n18311), .B2(n564), .ZN(n18691) );
  AOI22_X1 U10603 ( .A1(net716461), .A2(n568), .B1(n18347), .B2(n574), .ZN(
        n18680) );
  NOR2_X1 U10601 ( .A1(n588), .A2(net767232), .ZN(n18683) );
  OAI22_X1 U10600 ( .A1(n587), .A2(net767237), .B1(net716477), .B2(n24647), 
        .ZN(n18684) );
  AOI211_X1 U10599 ( .C1(n563), .C2(n18343), .A(n18683), .B(n18684), .ZN(
        n18682) );
  AOI22_X1 U10602 ( .A1(n18338), .A2(n572), .B1(n18339), .B2(n569), .ZN(n18681) );
  AOI22_X1 U10616 ( .A1(n18330), .A2(n570), .B1(n18331), .B2(n17716), .ZN(
        n18696) );
  AOI22_X1 U10614 ( .A1(n18325), .A2(n565), .B1(net716417), .B2(n24760), .ZN(
        n18698) );
  AOI22_X1 U10613 ( .A1(n18300), .A2(n566), .B1(net767235), .B2(n24761), .ZN(
        n18690) );
  AOI22_X1 U10615 ( .A1(net716423), .A2(n17715), .B1(net767214), .B2(n17717), 
        .ZN(n18697) );
  OAI22_X1 U10851 ( .A1(n708), .A2(n18315), .B1(n707), .B2(n18316), .ZN(n18987) );
  AOI22_X1 U10850 ( .A1(net767173), .A2(n691), .B1(n18321), .B2(n693), .ZN(
        n18989) );
  NAND2_X1 U10849 ( .A1(n18529), .A2(n685), .ZN(n18990) );
  OAI211_X1 U10848 ( .C1(n700), .C2(net518461), .A(n18989), .B(n18990), .ZN(
        n18988) );
  AOI211_X1 U10847 ( .C1(n18312), .C2(n694), .A(n18987), .B(n18988), .ZN(
        n18980) );
  AOI22_X1 U10853 ( .A1(n18307), .A2(n17741), .B1(net716405), .B2(n17740), 
        .ZN(n18994) );
  AOI22_X1 U10854 ( .A1(net767239), .A2(n24716), .B1(n18306), .B2(n695), .ZN(
        n18993) );
  AOI22_X1 U10855 ( .A1(n18310), .A2(n696), .B1(n18311), .B2(n682), .ZN(n18992) );
  AOI22_X1 U10846 ( .A1(net716461), .A2(n686), .B1(n18347), .B2(n692), .ZN(
        n18981) );
  NOR2_X1 U10844 ( .A1(n706), .A2(net767232), .ZN(n18984) );
  OAI22_X1 U10843 ( .A1(n705), .A2(net767237), .B1(net716477), .B2(n24642), 
        .ZN(n18985) );
  AOI211_X1 U10842 ( .C1(n681), .C2(n18343), .A(n18984), .B(n18985), .ZN(
        n18983) );
  AOI22_X1 U10845 ( .A1(n18338), .A2(n690), .B1(n18339), .B2(n687), .ZN(n18982) );
  AOI22_X1 U10859 ( .A1(n18330), .A2(n688), .B1(n18331), .B2(n17738), .ZN(
        n18997) );
  AOI22_X1 U10857 ( .A1(net767167), .A2(n683), .B1(n18326), .B2(n24750), .ZN(
        n18999) );
  AOI22_X1 U10856 ( .A1(n18300), .A2(n684), .B1(net767235), .B2(n24751), .ZN(
        n18991) );
  AOI22_X1 U10858 ( .A1(n18328), .A2(n17737), .B1(n18329), .B2(n17739), .ZN(
        n18998) );
  OAI22_X1 U10674 ( .A1(n669), .A2(n18315), .B1(n668), .B2(n18316), .ZN(n18767) );
  AOI22_X1 U10673 ( .A1(net767173), .A2(n652), .B1(n18321), .B2(n654), .ZN(
        n18769) );
  NAND2_X1 U10672 ( .A1(n18529), .A2(n646), .ZN(n18770) );
  OAI211_X1 U10671 ( .C1(n661), .C2(net518461), .A(n18769), .B(n18770), .ZN(
        n18768) );
  AOI211_X1 U10670 ( .C1(n18312), .C2(n655), .A(n18767), .B(n18768), .ZN(
        n18760) );
  AOI22_X1 U10676 ( .A1(n18307), .A2(n17734), .B1(net716405), .B2(n17733), 
        .ZN(n18774) );
  AOI22_X1 U10677 ( .A1(net767239), .A2(n24719), .B1(n18306), .B2(n656), .ZN(
        n18773) );
  AOI22_X1 U10678 ( .A1(n18310), .A2(n657), .B1(n18311), .B2(n643), .ZN(n18772) );
  AOI22_X1 U10669 ( .A1(net716461), .A2(n647), .B1(n18347), .B2(n653), .ZN(
        n18761) );
  NOR2_X1 U10667 ( .A1(n667), .A2(net767232), .ZN(n18764) );
  OAI22_X1 U10666 ( .A1(n666), .A2(net767237), .B1(net716477), .B2(n24645), 
        .ZN(n18765) );
  AOI211_X1 U10665 ( .C1(n642), .C2(n18343), .A(n18764), .B(n18765), .ZN(
        n18763) );
  AOI22_X1 U10668 ( .A1(n18338), .A2(n651), .B1(n18339), .B2(n648), .ZN(n18762) );
  AOI22_X1 U10682 ( .A1(n18330), .A2(n649), .B1(n18331), .B2(n17731), .ZN(
        n18777) );
  AOI22_X1 U10680 ( .A1(net767167), .A2(n644), .B1(n18326), .B2(n24756), .ZN(
        n18779) );
  AOI22_X1 U10679 ( .A1(n18300), .A2(n645), .B1(net767235), .B2(n24757), .ZN(
        n18771) );
  AOI22_X1 U10681 ( .A1(n18328), .A2(n17730), .B1(n18329), .B2(n17732), .ZN(
        n18778) );
  OAI22_X1 U10560 ( .A1(n437), .A2(n18315), .B1(n436), .B2(n18316), .ZN(n18632) );
  AOI22_X1 U10559 ( .A1(net767173), .A2(n420), .B1(n18321), .B2(n422), .ZN(
        n18634) );
  NAND2_X1 U10558 ( .A1(n18529), .A2(n414), .ZN(n18635) );
  OAI211_X1 U10557 ( .C1(n429), .C2(net518461), .A(n18634), .B(n18635), .ZN(
        n18633) );
  AOI211_X1 U10556 ( .C1(n18312), .C2(n423), .A(n18632), .B(n18633), .ZN(
        n18625) );
  AOI22_X1 U10562 ( .A1(n18307), .A2(n17694), .B1(net716405), .B2(n17693), 
        .ZN(n18639) );
  AOI22_X1 U10563 ( .A1(net767239), .A2(n24694), .B1(n18306), .B2(n424), .ZN(
        n18638) );
  AOI22_X1 U10564 ( .A1(n18310), .A2(n425), .B1(n18311), .B2(n411), .ZN(n18637) );
  AOI22_X1 U10555 ( .A1(net716461), .A2(n415), .B1(n18347), .B2(n421), .ZN(
        n18626) );
  NOR2_X1 U10553 ( .A1(n435), .A2(net767232), .ZN(n18629) );
  OAI22_X1 U10552 ( .A1(n434), .A2(net767237), .B1(net716477), .B2(n24626), 
        .ZN(n18630) );
  AOI211_X1 U10551 ( .C1(n410), .C2(n18343), .A(n18629), .B(n18630), .ZN(
        n18628) );
  AOI22_X1 U10554 ( .A1(n18338), .A2(n419), .B1(n18339), .B2(n416), .ZN(n18627) );
  AOI22_X1 U10572 ( .A1(n18330), .A2(n417), .B1(n18331), .B2(n17691), .ZN(
        n18642) );
  AOI22_X1 U10566 ( .A1(n18325), .A2(n412), .B1(net716417), .B2(n24745), .ZN(
        n18644) );
  AOI22_X1 U10565 ( .A1(n18300), .A2(n413), .B1(net767235), .B2(n24746), .ZN(
        n18636) );
  AOI22_X1 U10567 ( .A1(net716423), .A2(n17690), .B1(net767214), .B2(n17692), 
        .ZN(n18643) );
  AOI22_X1 U10837 ( .A1(n18330), .A2(n921), .B1(n18331), .B2(n17780), .ZN(
        n18970) );
  AOI22_X1 U10835 ( .A1(net767167), .A2(n916), .B1(net716417), .B2(n24739), 
        .ZN(n18972) );
  AOI22_X1 U10834 ( .A1(n18300), .A2(n917), .B1(net767235), .B2(n24740), .ZN(
        n18964) );
  AOI22_X1 U10836 ( .A1(n18328), .A2(n17779), .B1(n18329), .B2(n17781), .ZN(
        n18971) );
  OAI22_X1 U10740 ( .A1(n746), .A2(n18315), .B1(n745), .B2(n18316), .ZN(n18848) );
  AOI22_X1 U10739 ( .A1(net767173), .A2(n729), .B1(n18321), .B2(n731), .ZN(
        n18850) );
  NAND2_X1 U10738 ( .A1(n18529), .A2(n723), .ZN(n18851) );
  OAI211_X1 U10737 ( .C1(n738), .C2(net518461), .A(n18850), .B(n18851), .ZN(
        n18849) );
  AOI211_X1 U10736 ( .C1(n18312), .C2(n732), .A(n18848), .B(n18849), .ZN(
        n18841) );
  AOI22_X1 U10742 ( .A1(n18307), .A2(n17749), .B1(net716405), .B2(n17748), 
        .ZN(n18855) );
  AOI22_X1 U10743 ( .A1(net767239), .A2(n24692), .B1(n18306), .B2(n733), .ZN(
        n18854) );
  AOI22_X1 U10744 ( .A1(n18310), .A2(n734), .B1(n18311), .B2(n720), .ZN(n18853) );
  AOI22_X1 U10735 ( .A1(net716461), .A2(n724), .B1(n18347), .B2(n730), .ZN(
        n18842) );
  NOR2_X1 U10733 ( .A1(n744), .A2(net767232), .ZN(n18845) );
  OAI22_X1 U10732 ( .A1(n743), .A2(net767237), .B1(net716477), .B2(n24624), 
        .ZN(n18846) );
  AOI211_X1 U10731 ( .C1(n719), .C2(n18343), .A(n18845), .B(n18846), .ZN(
        n18844) );
  AOI22_X1 U10734 ( .A1(n18338), .A2(n728), .B1(n18339), .B2(n725), .ZN(n18843) );
  AOI22_X1 U10748 ( .A1(n18330), .A2(n726), .B1(n18331), .B2(n17746), .ZN(
        n18858) );
  AOI22_X1 U10746 ( .A1(net767167), .A2(n721), .B1(net716417), .B2(n24741), 
        .ZN(n18860) );
  AOI22_X1 U10745 ( .A1(n18300), .A2(n722), .B1(net767235), .B2(n24742), .ZN(
        n18852) );
  AOI22_X1 U10747 ( .A1(n18328), .A2(n17745), .B1(n18329), .B2(n17747), .ZN(
        n18859) );
  OAI22_X1 U10904 ( .A1(n2883), .A2(n18346), .B1(n2882), .B2(net767172), .ZN(
        n19041) );
  OAI22_X1 U10903 ( .A1(n2873), .A2(n18401), .B1(net767232), .B2(n24639), .ZN(
        n19042) );
  OAI22_X1 U10902 ( .A1(n2880), .A2(net716477), .B1(net767237), .B2(n24640), 
        .ZN(n19043) );
  OAI22_X1 U10901 ( .A1(n2879), .A2(n18369), .B1(n2877), .B2(n18361), .ZN(
        n19044) );
  NOR4_X1 U10900 ( .A1(n19041), .A2(n19042), .A3(n19043), .A4(n19044), .ZN(
        n19034) );
  AOI22_X1 U10899 ( .A1(n18300), .A2(n24714), .B1(net767235), .B2(n17822), 
        .ZN(n19035) );
  NOR2_X1 U10897 ( .A1(n2892), .A2(n18394), .ZN(n19038) );
  OAI22_X1 U10896 ( .A1(n2896), .A2(n18382), .B1(n2895), .B2(n18393), .ZN(
        n19039) );
  AOI211_X1 U10895 ( .C1(n17810), .C2(net767239), .A(n19038), .B(n19039), .ZN(
        n19037) );
  AOI22_X1 U10898 ( .A1(n18307), .A2(n17823), .B1(net716405), .B2(n17821), 
        .ZN(n19036) );
  AOI22_X1 U10906 ( .A1(net767167), .A2(n24713), .B1(n18326), .B2(n17811), 
        .ZN(n19050) );
  AOI22_X1 U10907 ( .A1(net767238), .A2(n17809), .B1(net767171), .B2(n17815), 
        .ZN(n19049) );
  AOI22_X1 U10908 ( .A1(net716423), .A2(n17813), .B1(net767214), .B2(n17816), 
        .ZN(n19048) );
  AOI22_X1 U10911 ( .A1(n18372), .A2(n17820), .B1(n18373), .B2(n17819), .ZN(
        n19054) );
  AOI22_X1 U10909 ( .A1(n18330), .A2(n24712), .B1(n18331), .B2(n17814), .ZN(
        n19047) );
  AOI22_X1 U11628 ( .A1(n19336), .A2(n843), .B1(n19337), .B2(n17766), .ZN(
        n19777) );
  AOI22_X1 U11625 ( .A1(n24026), .A2(n838), .B1(n19333), .B2(net741389), .ZN(
        n19779) );
  AOI22_X1 U11623 ( .A1(n19308), .A2(n839), .B1(n23995), .B2(net741388), .ZN(
        n19773) );
  AOI22_X1 U11627 ( .A1(n24007), .A2(n17765), .B1(n19335), .B2(n17767), .ZN(
        n19778) );
  AOI22_X1 U11619 ( .A1(n19315), .A2(n17769), .B1(n25683), .B2(n17768), .ZN(
        n19776) );
  AOI22_X1 U11620 ( .A1(n23994), .A2(net741442), .B1(n19314), .B2(n850), .ZN(
        n19775) );
  AOI22_X1 U11622 ( .A1(n19318), .A2(n851), .B1(n19319), .B2(n837), .ZN(n19774) );
  OAI22_X1 U11040 ( .A1(n2703), .A2(n18346), .B1(n2702), .B2(net767172), .ZN(
        n19208) );
  OAI22_X1 U11039 ( .A1(n2693), .A2(n18401), .B1(n18367), .B2(n24629), .ZN(
        n19209) );
  OAI22_X1 U11038 ( .A1(n2700), .A2(net716477), .B1(net767237), .B2(n24630), 
        .ZN(n19210) );
  OAI22_X1 U11037 ( .A1(n2699), .A2(n18369), .B1(n2697), .B2(n18361), .ZN(
        n19211) );
  NOR4_X1 U11036 ( .A1(n19208), .A2(n19209), .A3(n19210), .A4(n19211), .ZN(
        n19201) );
  AOI22_X1 U11035 ( .A1(n18300), .A2(n24700), .B1(net767235), .B2(n18017), 
        .ZN(n19202) );
  NOR2_X1 U11033 ( .A1(n2712), .A2(n18394), .ZN(n19205) );
  OAI22_X1 U11032 ( .A1(n2716), .A2(n18382), .B1(n2715), .B2(n18393), .ZN(
        n19206) );
  AOI211_X1 U11031 ( .C1(n18005), .C2(net767239), .A(n19205), .B(n19206), .ZN(
        n19204) );
  AOI22_X1 U11034 ( .A1(n18307), .A2(n18018), .B1(net716405), .B2(n18016), 
        .ZN(n19203) );
  AOI22_X1 U11042 ( .A1(net767167), .A2(n24699), .B1(net716417), .B2(n18006), 
        .ZN(n19217) );
  AOI22_X1 U11043 ( .A1(net767238), .A2(n18004), .B1(net767171), .B2(n18010), 
        .ZN(n19216) );
  AOI22_X1 U11044 ( .A1(net716423), .A2(n18008), .B1(net767214), .B2(n18011), 
        .ZN(n19215) );
  AOI22_X1 U11047 ( .A1(n18372), .A2(n18015), .B1(n18373), .B2(n18014), .ZN(
        n19221) );
  AOI22_X1 U11045 ( .A1(n18330), .A2(n24698), .B1(n18331), .B2(n18009), .ZN(
        n19214) );
  OAI22_X1 U11392 ( .A1(n437), .A2(n19323), .B1(n436), .B2(n19324), .ZN(n19571) );
  AOI22_X1 U11391 ( .A1(n19327), .A2(n420), .B1(n19328), .B2(n422), .ZN(n19573) );
  NAND2_X1 U11390 ( .A1(n19530), .A2(n414), .ZN(n19574) );
  OAI211_X1 U11389 ( .C1(n429), .C2(n26785), .A(n19573), .B(n19574), .ZN(
        n19572) );
  AOI211_X1 U11388 ( .C1(n19320), .C2(n423), .A(n19571), .B(n19572), .ZN(
        n19565) );
  AOI22_X1 U11387 ( .A1(n25679), .A2(n415), .B1(n25666), .B2(n421), .ZN(n19566) );
  NOR2_X1 U11385 ( .A1(n435), .A2(n25677), .ZN(n19569) );
  OAI22_X1 U11384 ( .A1(n434), .A2(n25675), .B1(n25678), .B2(n24626), .ZN(
        n19570) );
  AOI211_X1 U11383 ( .C1(n410), .C2(n19348), .A(n19569), .B(n19570), .ZN(
        n19568) );
  AOI22_X1 U11386 ( .A1(n19344), .A2(n419), .B1(n19345), .B2(n416), .ZN(n19567) );
  AOI22_X1 U11403 ( .A1(n19336), .A2(n417), .B1(n19337), .B2(n17691), .ZN(
        n19579) );
  AOI22_X1 U11400 ( .A1(n24026), .A2(n412), .B1(n25682), .B2(n24745), .ZN(
        n19581) );
  AOI22_X1 U11398 ( .A1(n19308), .A2(n413), .B1(n23995), .B2(n24746), .ZN(
        n19575) );
  AOI22_X1 U11402 ( .A1(n19334), .A2(n17690), .B1(n25681), .B2(n17692), .ZN(
        n19580) );
  AOI22_X1 U11394 ( .A1(n19315), .A2(n17694), .B1(n25683), .B2(n17693), .ZN(
        n19578) );
  AOI22_X1 U11395 ( .A1(n23994), .A2(n24694), .B1(n19314), .B2(n424), .ZN(
        n19577) );
  AOI22_X1 U11397 ( .A1(n19318), .A2(n425), .B1(n19319), .B2(n411), .ZN(n19576) );
  OAI22_X1 U11517 ( .A1(n669), .A2(n19323), .B1(n668), .B2(n19324), .ZN(n19681) );
  AOI22_X1 U11516 ( .A1(n19327), .A2(n652), .B1(n19328), .B2(n654), .ZN(n19683) );
  NAND2_X1 U11515 ( .A1(n19530), .A2(n646), .ZN(n19684) );
  OAI211_X1 U11514 ( .C1(n661), .C2(n26785), .A(n19683), .B(n19684), .ZN(
        n19682) );
  AOI211_X1 U11513 ( .C1(n19320), .C2(n655), .A(n19681), .B(n19682), .ZN(
        n19675) );
  AOI22_X1 U11512 ( .A1(n25679), .A2(n647), .B1(n25666), .B2(n653), .ZN(n19676) );
  NOR2_X1 U11510 ( .A1(n667), .A2(n25677), .ZN(n19679) );
  OAI22_X1 U11509 ( .A1(n666), .A2(n25676), .B1(n25678), .B2(n24645), .ZN(
        n19680) );
  AOI211_X1 U11508 ( .C1(n642), .C2(n19348), .A(n19679), .B(n19680), .ZN(
        n19678) );
  AOI22_X1 U11511 ( .A1(n19344), .A2(n651), .B1(n19345), .B2(n648), .ZN(n19677) );
  AOI22_X1 U11528 ( .A1(n19336), .A2(n649), .B1(n19337), .B2(n17731), .ZN(
        n19689) );
  AOI22_X1 U11525 ( .A1(n24026), .A2(n644), .B1(n19333), .B2(n24756), .ZN(
        n19691) );
  AOI22_X1 U11523 ( .A1(n19308), .A2(n645), .B1(n23995), .B2(n24757), .ZN(
        n19685) );
  AOI22_X1 U11527 ( .A1(n24007), .A2(n17730), .B1(n25681), .B2(n17732), .ZN(
        n19690) );
  AOI22_X1 U11519 ( .A1(n19315), .A2(n17734), .B1(n25683), .B2(n17733), .ZN(
        n19688) );
  AOI22_X1 U11520 ( .A1(n23994), .A2(n24719), .B1(n19314), .B2(n656), .ZN(
        n19687) );
  AOI22_X1 U11522 ( .A1(n19318), .A2(n657), .B1(n19319), .B2(n643), .ZN(n19686) );
  AOI22_X1 U11914 ( .A1(n24026), .A2(n24702), .B1(n19333), .B2(n17879), .ZN(
        n20013) );
  AOI22_X1 U11916 ( .A1(n25674), .A2(n17877), .B1(n25680), .B2(n17883), .ZN(
        n20012) );
  AOI22_X1 U11917 ( .A1(n24007), .A2(n17881), .B1(n19335), .B2(n17884), .ZN(
        n20011) );
  OAI22_X1 U11694 ( .A1(n941), .A2(n19323), .B1(n940), .B2(n19324), .ZN(n19835) );
  AOI22_X1 U11693 ( .A1(n19327), .A2(n924), .B1(n19328), .B2(n926), .ZN(n19837) );
  NAND2_X1 U11692 ( .A1(n19530), .A2(n918), .ZN(n19838) );
  OAI211_X1 U11691 ( .C1(n933), .C2(n26785), .A(n19837), .B(n19838), .ZN(
        n19836) );
  AOI211_X1 U11690 ( .C1(n19320), .C2(n927), .A(n19835), .B(n19836), .ZN(
        n19829) );
  AOI22_X1 U11689 ( .A1(n25679), .A2(n919), .B1(n25667), .B2(n925), .ZN(n19830) );
  NOR2_X1 U11687 ( .A1(n939), .A2(n25677), .ZN(n19833) );
  OAI22_X1 U11686 ( .A1(n938), .A2(n25675), .B1(n25678), .B2(n24622), .ZN(
        n19834) );
  AOI211_X1 U11685 ( .C1(n914), .C2(n19348), .A(n19833), .B(n19834), .ZN(
        n19832) );
  AOI22_X1 U11688 ( .A1(n19344), .A2(n923), .B1(n19345), .B2(n920), .ZN(n19831) );
  AOI22_X1 U11705 ( .A1(n19336), .A2(n921), .B1(n19337), .B2(n17780), .ZN(
        n19843) );
  AOI22_X1 U11702 ( .A1(n24026), .A2(n916), .B1(n19333), .B2(n24739), .ZN(
        n19845) );
  AOI22_X1 U11700 ( .A1(n19308), .A2(n917), .B1(n23995), .B2(n24740), .ZN(
        n19839) );
  AOI22_X1 U11704 ( .A1(n24007), .A2(n17779), .B1(n25681), .B2(n17781), .ZN(
        n19844) );
  AOI22_X1 U11696 ( .A1(n19315), .A2(n17783), .B1(n25683), .B2(n17782), .ZN(
        n19842) );
  AOI22_X1 U11697 ( .A1(n23994), .A2(n24691), .B1(n19314), .B2(n928), .ZN(
        n19841) );
  AOI22_X1 U11699 ( .A1(n19318), .A2(n929), .B1(n19319), .B2(n915), .ZN(n19840) );
  OAI22_X1 U11492 ( .A1(n399), .A2(n19323), .B1(n398), .B2(n19324), .ZN(n19659) );
  AOI22_X1 U11491 ( .A1(n19327), .A2(n382), .B1(n19328), .B2(n384), .ZN(n19661) );
  NAND2_X1 U11490 ( .A1(n19530), .A2(n376), .ZN(n19662) );
  OAI211_X1 U11489 ( .C1(n391), .C2(n26785), .A(n19661), .B(n19662), .ZN(
        n19660) );
  AOI211_X1 U11488 ( .C1(n19320), .C2(n385), .A(n19659), .B(n19660), .ZN(
        n19653) );
  AOI22_X1 U11487 ( .A1(n25679), .A2(n377), .B1(n25666), .B2(n383), .ZN(n19654) );
  NOR2_X1 U11485 ( .A1(n397), .A2(n25677), .ZN(n19657) );
  OAI22_X1 U11484 ( .A1(n396), .A2(n25676), .B1(n25678), .B2(n24646), .ZN(
        n19658) );
  AOI211_X1 U11483 ( .C1(n372), .C2(n19348), .A(n19657), .B(n19658), .ZN(
        n19656) );
  AOI22_X1 U11486 ( .A1(n19344), .A2(n381), .B1(n19345), .B2(n378), .ZN(n19655) );
  AOI22_X1 U11503 ( .A1(n19336), .A2(n379), .B1(n19337), .B2(n17684), .ZN(
        n19667) );
  AOI22_X1 U11500 ( .A1(n24026), .A2(n374), .B1(n25682), .B2(n24758), .ZN(
        n19669) );
  AOI22_X1 U11498 ( .A1(n19308), .A2(n375), .B1(n23995), .B2(n24759), .ZN(
        n19663) );
  AOI22_X1 U11502 ( .A1(n24007), .A2(n17683), .B1(n19335), .B2(n17685), .ZN(
        n19668) );
  AOI22_X1 U11494 ( .A1(n19315), .A2(n17687), .B1(n25683), .B2(n17686), .ZN(
        n19666) );
  AOI22_X1 U11495 ( .A1(n23994), .A2(n24720), .B1(n19314), .B2(n386), .ZN(
        n19665) );
  AOI22_X1 U11497 ( .A1(n19318), .A2(n387), .B1(n19319), .B2(n373), .ZN(n19664) );
  OAI22_X1 U11567 ( .A1(n823), .A2(n19323), .B1(n822), .B2(n19324), .ZN(n19725) );
  AOI22_X1 U11566 ( .A1(n19327), .A2(n806), .B1(n19328), .B2(n808), .ZN(n19727) );
  NAND2_X1 U11565 ( .A1(n19530), .A2(n800), .ZN(n19728) );
  OAI211_X1 U11564 ( .C1(n815), .C2(n26785), .A(n19727), .B(n19728), .ZN(
        n19726) );
  AOI211_X1 U11563 ( .C1(n19320), .C2(n809), .A(n19725), .B(n19726), .ZN(
        n19719) );
  AOI22_X1 U11562 ( .A1(n25679), .A2(n801), .B1(n19351), .B2(n807), .ZN(n19720) );
  NOR2_X1 U11560 ( .A1(n821), .A2(n25677), .ZN(n19723) );
  OAI22_X1 U11559 ( .A1(n820), .A2(n25675), .B1(n25678), .B2(net741518), .ZN(
        n19724) );
  AOI211_X1 U11558 ( .C1(n796), .C2(n19348), .A(n19723), .B(n19724), .ZN(
        n19722) );
  AOI22_X1 U11561 ( .A1(n19344), .A2(n805), .B1(n19345), .B2(n802), .ZN(n19721) );
  AOI22_X1 U11578 ( .A1(n19336), .A2(n803), .B1(n19337), .B2(n17759), .ZN(
        n19733) );
  AOI22_X1 U11575 ( .A1(n24026), .A2(n798), .B1(n19333), .B2(net741385), .ZN(
        n19735) );
  AOI22_X1 U11573 ( .A1(n19308), .A2(n799), .B1(n23995), .B2(net741384), .ZN(
        n19729) );
  AOI22_X1 U11577 ( .A1(n24007), .A2(n17758), .B1(n19335), .B2(n17760), .ZN(
        n19734) );
  AOI22_X1 U11569 ( .A1(n19315), .A2(n17762), .B1(n25683), .B2(n17761), .ZN(
        n19732) );
  AOI22_X1 U11570 ( .A1(n23994), .A2(net741440), .B1(n19314), .B2(n810), .ZN(
        n19731) );
  AOI22_X1 U11572 ( .A1(n19318), .A2(n811), .B1(n19319), .B2(n797), .ZN(n19730) );
  OAI22_X1 U11542 ( .A1(n784), .A2(n19323), .B1(n783), .B2(n19324), .ZN(n19703) );
  AOI22_X1 U11541 ( .A1(n19327), .A2(n767), .B1(n19328), .B2(n769), .ZN(n19705) );
  NAND2_X1 U11540 ( .A1(n19530), .A2(n761), .ZN(n19706) );
  OAI211_X1 U11539 ( .C1(n776), .C2(n26785), .A(n19705), .B(n19706), .ZN(
        n19704) );
  AOI211_X1 U11538 ( .C1(n19320), .C2(n770), .A(n19703), .B(n19704), .ZN(
        n19697) );
  AOI22_X1 U11537 ( .A1(n25679), .A2(n762), .B1(n19351), .B2(n768), .ZN(n19698) );
  NOR2_X1 U11535 ( .A1(n782), .A2(n25677), .ZN(n19701) );
  OAI22_X1 U11534 ( .A1(n781), .A2(n25675), .B1(n25678), .B2(n24644), .ZN(
        n19702) );
  AOI211_X1 U11533 ( .C1(n757), .C2(n19348), .A(n19701), .B(n19702), .ZN(
        n19700) );
  AOI22_X1 U11536 ( .A1(n19344), .A2(n766), .B1(n19345), .B2(n763), .ZN(n19699) );
  AOI22_X1 U11553 ( .A1(n19336), .A2(n764), .B1(n19337), .B2(n17752), .ZN(
        n19711) );
  AOI22_X1 U11550 ( .A1(n24026), .A2(n759), .B1(n19333), .B2(n24754), .ZN(
        n19713) );
  AOI22_X1 U11548 ( .A1(n19308), .A2(n760), .B1(n23995), .B2(n24755), .ZN(
        n19707) );
  AOI22_X1 U11552 ( .A1(n24007), .A2(n17751), .B1(n25681), .B2(n17753), .ZN(
        n19712) );
  AOI22_X1 U11544 ( .A1(n19315), .A2(n17755), .B1(n25683), .B2(n17754), .ZN(
        n19710) );
  AOI22_X1 U11545 ( .A1(n23994), .A2(n24718), .B1(n19314), .B2(n771), .ZN(
        n19709) );
  AOI22_X1 U11547 ( .A1(n19318), .A2(n772), .B1(n19319), .B2(n758), .ZN(n19708) );
  OAI22_X1 U10974 ( .A1(n2991), .A2(n18346), .B1(n2990), .B2(net767172), .ZN(
        n19124) );
  OAI22_X1 U10973 ( .A1(n2981), .A2(n18401), .B1(net767232), .B2(n24620), .ZN(
        n19125) );
  OAI22_X1 U10972 ( .A1(n2988), .A2(net716477), .B1(net767237), .B2(n24621), 
        .ZN(n19126) );
  OAI22_X1 U10971 ( .A1(n2987), .A2(n18369), .B1(n2985), .B2(n18361), .ZN(
        n19127) );
  NOR4_X1 U10970 ( .A1(n19124), .A2(n19125), .A3(n19126), .A4(n19127), .ZN(
        n19117) );
  AOI22_X1 U10969 ( .A1(n18300), .A2(n24684), .B1(net767235), .B2(n17856), 
        .ZN(n19118) );
  NOR2_X1 U10967 ( .A1(n3000), .A2(n18394), .ZN(n19121) );
  OAI22_X1 U10966 ( .A1(n3004), .A2(n18382), .B1(n3003), .B2(n18393), .ZN(
        n19122) );
  AOI211_X1 U10965 ( .C1(n17844), .C2(net767239), .A(n19121), .B(n19122), .ZN(
        n19120) );
  AOI22_X1 U10968 ( .A1(n18307), .A2(n17857), .B1(net716405), .B2(n17855), 
        .ZN(n19119) );
  AOI22_X1 U10976 ( .A1(net767167), .A2(n24683), .B1(n18326), .B2(n17845), 
        .ZN(n19133) );
  AOI22_X1 U10977 ( .A1(net767238), .A2(n17843), .B1(net767171), .B2(n17849), 
        .ZN(n19132) );
  AOI22_X1 U10978 ( .A1(net716423), .A2(n17847), .B1(net767214), .B2(n17850), 
        .ZN(n19131) );
  AOI22_X1 U10981 ( .A1(n18372), .A2(n17854), .B1(n18373), .B2(n17853), .ZN(
        n19137) );
  AOI22_X1 U10979 ( .A1(n18330), .A2(n24682), .B1(n18331), .B2(n17848), .ZN(
        n19130) );
  NOR2_X1 U10346 ( .A1(n363), .A2(net741544), .ZN(n18301) );
  AOI22_X1 U10345 ( .A1(n18307), .A2(n17681), .B1(net716405), .B2(n17680), 
        .ZN(n18304) );
  NAND2_X1 U10344 ( .A1(n18306), .A2(n348), .ZN(n18305) );
  OAI211_X1 U10343 ( .C1(n351), .C2(net741541), .A(n18304), .B(n18305), .ZN(
        n18302) );
  AOI211_X1 U10342 ( .C1(n337), .C2(n18300), .A(n18301), .B(n18302), .ZN(
        n18299) );
  AOI22_X1 U10351 ( .A1(net767173), .A2(n344), .B1(n18321), .B2(n346), .ZN(
        n18296) );
  OAI22_X1 U10350 ( .A1(n353), .A2(net518461), .B1(n18318), .B2(n24667), .ZN(
        n18313) );
  OAI22_X1 U10349 ( .A1(n361), .A2(n18315), .B1(n360), .B2(n18316), .ZN(n18314) );
  AOI211_X1 U10348 ( .C1(n18312), .C2(n347), .A(n18313), .B(n18314), .ZN(
        n18297) );
  AOI22_X1 U10347 ( .A1(n18310), .A2(n349), .B1(n18311), .B2(n335), .ZN(n18298) );
  AOI22_X1 U10360 ( .A1(net716461), .A2(n339), .B1(n18347), .B2(n345), .ZN(
        n18334) );
  AOI22_X1 U10358 ( .A1(net741539), .A2(n342), .B1(net741532), .B2(n24771), 
        .ZN(n18336) );
  AOI22_X1 U10357 ( .A1(n18338), .A2(n343), .B1(n18339), .B2(n340), .ZN(n18337) );
  AOI22_X1 U10359 ( .A1(n18343), .A2(n334), .B1(net716491), .B2(n24770), .ZN(
        n18335) );
  AOI22_X1 U10352 ( .A1(net767167), .A2(n336), .B1(net716417), .B2(n24772), 
        .ZN(n18324) );
  AOI22_X1 U10353 ( .A1(n18328), .A2(n17677), .B1(net767214), .B2(n17679), 
        .ZN(n18323) );
  AOI22_X1 U10354 ( .A1(n18330), .A2(n341), .B1(n18331), .B2(n17678), .ZN(
        n18322) );
  OAI22_X1 U11312 ( .A1(n465), .A2(n26785), .B1(n19326), .B2(n24654), .ZN(
        n19506) );
  OAI22_X1 U11311 ( .A1(n473), .A2(n19323), .B1(n472), .B2(n19324), .ZN(n19507) );
  AOI211_X1 U11310 ( .C1(n19320), .C2(n459), .A(n19506), .B(n19507), .ZN(
        n19500) );
  OAI22_X1 U11307 ( .A1(n474), .A2(n24613), .B1(n19390), .B2(n24655), .ZN(
        n19503) );
  OAI22_X1 U11305 ( .A1(n463), .A2(n24614), .B1(n19389), .B2(n24656), .ZN(
        n19504) );
  OAI22_X1 U11303 ( .A1(n1755), .A2(n24615), .B1(n475), .B2(n19384), .ZN(
        n19505) );
  NOR3_X1 U11302 ( .A1(n19503), .A2(n19504), .A3(n19505), .ZN(n19502) );
  AOI22_X1 U11313 ( .A1(n19327), .A2(n456), .B1(n19328), .B2(n458), .ZN(n19499) );
  AOI22_X1 U11309 ( .A1(n19318), .A2(n461), .B1(n19319), .B2(n447), .ZN(n19501) );
  AOI22_X1 U11328 ( .A1(n25679), .A2(n451), .B1(n25667), .B2(n457), .ZN(n19511) );
  AOI22_X1 U11321 ( .A1(n19344), .A2(n455), .B1(n19345), .B2(n452), .ZN(n19514) );
  AOI22_X1 U11322 ( .A1(n24617), .A2(n454), .B1(n24591), .B2(n24767), .ZN(
        n19513) );
  AOI22_X1 U11326 ( .A1(n19348), .A2(n446), .B1(n24619), .B2(n24766), .ZN(
        n19512) );
  AOI22_X1 U11314 ( .A1(n24026), .A2(n448), .B1(n25682), .B2(n24769), .ZN(
        n19510) );
  AOI22_X1 U11316 ( .A1(n19334), .A2(n17697), .B1(n25681), .B2(n24768), .ZN(
        n19509) );
  AOI22_X1 U11318 ( .A1(n19336), .A2(n453), .B1(n19337), .B2(n17698), .ZN(
        n19508) );
  OAI22_X1 U11341 ( .A1(n511), .A2(n19323), .B1(n510), .B2(n19324), .ZN(n19526) );
  AOI22_X1 U11340 ( .A1(n19327), .A2(n494), .B1(n19328), .B2(n496), .ZN(n19528) );
  NAND2_X1 U11339 ( .A1(n19530), .A2(n488), .ZN(n19529) );
  OAI211_X1 U11338 ( .C1(n503), .C2(n26785), .A(n19528), .B(n19529), .ZN(
        n19527) );
  AOI211_X1 U11337 ( .C1(n19320), .C2(n497), .A(n19526), .B(n19527), .ZN(
        n19520) );
  AOI22_X1 U11336 ( .A1(n25679), .A2(n489), .B1(n25666), .B2(n495), .ZN(n19521) );
  NOR2_X1 U11334 ( .A1(n509), .A2(n25677), .ZN(n19524) );
  OAI22_X1 U11333 ( .A1(n508), .A2(n25675), .B1(n25678), .B2(n24653), .ZN(
        n19525) );
  AOI211_X1 U11332 ( .C1(n484), .C2(n19348), .A(n19524), .B(n19525), .ZN(
        n19523) );
  AOI22_X1 U11335 ( .A1(n19344), .A2(n493), .B1(n19345), .B2(n490), .ZN(n19522) );
  AOI22_X1 U11352 ( .A1(n19336), .A2(n491), .B1(n19337), .B2(n17702), .ZN(
        n19535) );
  AOI22_X1 U11349 ( .A1(n24026), .A2(n486), .B1(n25682), .B2(n24764), .ZN(
        n19537) );
  AOI22_X1 U11347 ( .A1(n19308), .A2(n487), .B1(n23995), .B2(n24765), .ZN(
        n19531) );
  AOI22_X1 U11351 ( .A1(n19334), .A2(n17701), .B1(n25681), .B2(n17703), .ZN(
        n19536) );
  AOI22_X1 U11343 ( .A1(n19315), .A2(n17705), .B1(n25683), .B2(n17704), .ZN(
        n19534) );
  AOI22_X1 U11344 ( .A1(n23994), .A2(n24723), .B1(n19314), .B2(n498), .ZN(
        n19533) );
  AOI22_X1 U11346 ( .A1(n19318), .A2(n499), .B1(n19319), .B2(n485), .ZN(n19532) );
  OAI22_X1 U10366 ( .A1(n18363), .A2(n24590), .B1(n18332), .B2(n24666), .ZN(
        n18359) );
  OAI22_X1 U10367 ( .A1(n2016), .A2(net716477), .B1(net767232), .B2(n24665), 
        .ZN(n18358) );
  OAI22_X1 U10365 ( .A1(n2013), .A2(n18361), .B1(n2012), .B2(n18362), .ZN(
        n18360) );
  OAI22_X1 U10379 ( .A1(n2031), .A2(n18393), .B1(n2028), .B2(n18394), .ZN(
        n18392) );
  AOI21_X1 U10378 ( .B1(net767239), .B2(n17895), .A(n18392), .ZN(n18383) );
  OAI22_X1 U10377 ( .A1(n2025), .A2(n18390), .B1(n2010), .B2(n18318), .ZN(
        n18385) );
  OAI22_X1 U10376 ( .A1(n2029), .A2(n18387), .B1(n18388), .B2(n24663), .ZN(
        n18386) );
  AOI211_X1 U10375 ( .C1(net716405), .C2(n17905), .A(n18385), .B(n18386), .ZN(
        n18384) );
  OAI211_X1 U10374 ( .C1(n2032), .C2(n18382), .A(n18383), .B(n18384), .ZN(
        n18381) );
  AOI22_X1 U10381 ( .A1(net716417), .A2(n17896), .B1(net767235), .B2(n17906), 
        .ZN(n18396) );
  OAI21_X1 U10380 ( .B1(n2034), .B2(n18395), .A(n18396), .ZN(n18380) );
  OAI22_X1 U10383 ( .A1(n2026), .A2(n18400), .B1(n2009), .B2(n18401), .ZN(
        n18399) );
  OAI22_X1 U10368 ( .A1(n2015), .A2(n18369), .B1(net767237), .B2(n24664), .ZN(
        n18357) );
  OAI22_X1 U11225 ( .A1(n19367), .A2(n24593), .B1(n19338), .B2(n24673), .ZN(
        n19429) );
  OAI22_X1 U11226 ( .A1(n2088), .A2(n25678), .B1(n25677), .B2(n24658), .ZN(
        n19428) );
  OAI22_X1 U11224 ( .A1(n2085), .A2(n19365), .B1(n2084), .B2(n19366), .ZN(
        n19430) );
  OAI22_X1 U11240 ( .A1(n2103), .A2(n19388), .B1(n2100), .B2(n19389), .ZN(
        n19439) );
  AOI21_X1 U11239 ( .B1(n23994), .B2(n17926), .A(n19439), .ZN(n19435) );
  OAI22_X1 U11238 ( .A1(n2097), .A2(n19385), .B1(n2082), .B2(n19326), .ZN(
        n19437) );
  OAI22_X1 U11237 ( .A1(n2101), .A2(n19383), .B1(n19384), .B2(n24671), .ZN(
        n19438) );
  AOI211_X1 U11236 ( .C1(n25683), .C2(n17936), .A(n19437), .B(n19438), .ZN(
        n19436) );
  OAI211_X1 U11235 ( .C1(n2104), .C2(n19378), .A(n19435), .B(n19436), .ZN(
        n19434) );
  AOI22_X1 U11242 ( .A1(n25682), .A2(n17927), .B1(n23995), .B2(n17937), .ZN(
        n19440) );
  OAI21_X1 U11241 ( .B1(n2106), .B2(n19390), .A(n19440), .ZN(n19433) );
  OAI22_X1 U11245 ( .A1(n2098), .A2(n19395), .B1(n2081), .B2(n19396), .ZN(
        n19441) );
  OAI22_X1 U11227 ( .A1(n2087), .A2(n19370), .B1(n25676), .B2(n24672), .ZN(
        n19427) );
  OAI22_X1 U10435 ( .A1(n24592), .A2(n18363), .B1(n24670), .B2(n18332), .ZN(
        n18476) );
  OAI22_X1 U10436 ( .A1(n2124), .A2(net716477), .B1(net767232), .B2(n24657), 
        .ZN(n18475) );
  OAI22_X1 U10434 ( .A1(n2120), .A2(n18362), .B1(n2121), .B2(n18361), .ZN(
        n18477) );
  OAI22_X1 U10448 ( .A1(n2136), .A2(n18394), .B1(n2139), .B2(n18393), .ZN(
        n18495) );
  AOI21_X1 U10447 ( .B1(n17942), .B2(net767239), .A(n18495), .ZN(n18490) );
  OAI22_X1 U10446 ( .A1(n2118), .A2(n18318), .B1(n2133), .B2(n18390), .ZN(
        n18492) );
  OAI22_X1 U10445 ( .A1(n2137), .A2(n18387), .B1(n24668), .B2(n18388), .ZN(
        n18493) );
  AOI211_X1 U10444 ( .C1(n17952), .C2(net716405), .A(n18492), .B(n18493), .ZN(
        n18491) );
  OAI211_X1 U10443 ( .C1(n2140), .C2(n18382), .A(n18490), .B(n18491), .ZN(
        n18489) );
  AOI22_X1 U10450 ( .A1(n17943), .A2(net716417), .B1(n17953), .B2(net767235), 
        .ZN(n18496) );
  OAI21_X1 U10449 ( .B1(n2142), .B2(n18395), .A(n18496), .ZN(n18488) );
  OAI22_X1 U10452 ( .A1(n2117), .A2(n18401), .B1(n2134), .B2(n18400), .ZN(
        n18497) );
  OAI22_X1 U10437 ( .A1(n2123), .A2(n18369), .B1(n24669), .B2(net767237), .ZN(
        n18474) );
  OAI22_X1 U11251 ( .A1(n19367), .A2(n24592), .B1(n19338), .B2(n24670), .ZN(
        n19451) );
  OAI22_X1 U11252 ( .A1(n2124), .A2(n25678), .B1(n25677), .B2(n24657), .ZN(
        n19450) );
  OAI22_X1 U11250 ( .A1(n2121), .A2(n19365), .B1(n2120), .B2(n19366), .ZN(
        n19452) );
  OAI22_X1 U11266 ( .A1(n2139), .A2(n19388), .B1(n2136), .B2(n19389), .ZN(
        n19461) );
  AOI21_X1 U11265 ( .B1(n23994), .B2(n17942), .A(n19461), .ZN(n19457) );
  OAI22_X1 U11264 ( .A1(n2133), .A2(n19385), .B1(n2118), .B2(n19326), .ZN(
        n19459) );
  OAI22_X1 U11263 ( .A1(n2137), .A2(n19383), .B1(n19384), .B2(n24668), .ZN(
        n19460) );
  AOI211_X1 U11262 ( .C1(n25683), .C2(n17952), .A(n19459), .B(n19460), .ZN(
        n19458) );
  OAI211_X1 U11261 ( .C1(n2140), .C2(n19378), .A(n19457), .B(n19458), .ZN(
        n19456) );
  AOI22_X1 U11268 ( .A1(n25682), .A2(n17943), .B1(n23995), .B2(n17953), .ZN(
        n19462) );
  OAI21_X1 U11267 ( .B1(n2142), .B2(n19390), .A(n19462), .ZN(n19455) );
  OAI22_X1 U11271 ( .A1(n2134), .A2(n19395), .B1(n2117), .B2(n19396), .ZN(
        n19463) );
  OAI22_X1 U11253 ( .A1(n2123), .A2(n19370), .B1(n25675), .B2(n24669), .ZN(
        n19449) );
  OAI22_X1 U11636 ( .A1(n24676), .A2(n19367), .B1(n24594), .B2(n19338), .ZN(
        n19789) );
  OAI22_X1 U11637 ( .A1(n2304), .A2(n25678), .B1(n25677), .B2(n24623), .ZN(
        n19788) );
  OAI22_X1 U11635 ( .A1(n2300), .A2(n19366), .B1(n2301), .B2(n19365), .ZN(
        n19790) );
  OAI22_X1 U11651 ( .A1(n2316), .A2(n19389), .B1(n2319), .B2(n19388), .ZN(
        n19799) );
  AOI21_X1 U11650 ( .B1(n17990), .B2(n23994), .A(n19799), .ZN(n19795) );
  OAI22_X1 U11649 ( .A1(n2298), .A2(n19326), .B1(n2313), .B2(n19385), .ZN(
        n19797) );
  OAI22_X1 U11648 ( .A1(n2317), .A2(n19383), .B1(n24674), .B2(n19384), .ZN(
        n19798) );
  AOI211_X1 U11647 ( .C1(n18000), .C2(n25683), .A(n19797), .B(n19798), .ZN(
        n19796) );
  OAI211_X1 U11646 ( .C1(n2320), .C2(n19378), .A(n19795), .B(n19796), .ZN(
        n19794) );
  AOI22_X1 U11653 ( .A1(n17991), .A2(n25682), .B1(n18001), .B2(n23995), .ZN(
        n19800) );
  OAI21_X1 U11652 ( .B1(n2322), .B2(n19390), .A(n19800), .ZN(n19793) );
  OAI22_X1 U11656 ( .A1(n2297), .A2(n19396), .B1(n2314), .B2(n19395), .ZN(
        n19801) );
  OAI22_X1 U11638 ( .A1(n2303), .A2(n19370), .B1(n24675), .B2(n25676), .ZN(
        n19787) );
  AOI22_X1 U11844 ( .A1(n19372), .A2(n17803), .B1(n19373), .B2(n17802), .ZN(
        n19952) );
  AOI22_X1 U11838 ( .A1(n24026), .A2(n995), .B1(n19333), .B2(n17795), .ZN(
        n19950) );
  AOI22_X1 U11841 ( .A1(n19336), .A2(n24707), .B1(n19337), .B2(n14402), .ZN(
        n19947) );
  AOI22_X1 U11840 ( .A1(n24007), .A2(n17797), .B1(n25681), .B2(n17799), .ZN(
        n19948) );
  AOI22_X1 U11839 ( .A1(n25674), .A2(n17793), .B1(n25680), .B2(n17798), .ZN(
        n19949) );
  AOI22_X1 U11830 ( .A1(n19308), .A2(n996), .B1(n23995), .B2(n17805), .ZN(
        n19941) );
  AOI22_X1 U11826 ( .A1(n19318), .A2(n24708), .B1(n19319), .B2(n994), .ZN(
        n19942) );
  AOI22_X1 U11823 ( .A1(n23994), .A2(n17794), .B1(n19314), .B2(n24747), .ZN(
        n19943) );
  AOI22_X1 U11822 ( .A1(n19315), .A2(n17806), .B1(n25683), .B2(n17804), .ZN(
        n19944) );
  NAND4_X1 U11821 ( .A1(n19941), .A2(n19942), .A3(n19943), .A4(n19944), .ZN(
        n19940) );
  OAI22_X1 U11835 ( .A1(n2951), .A2(n19370), .B1(n19365), .B2(n24636), .ZN(
        n19938) );
  AOI22_X1 U11833 ( .A1(n19348), .A2(n993), .B1(n24619), .B2(n17801), .ZN(
        n19945) );
  NAND2_X1 U11832 ( .A1(n25679), .A2(n998), .ZN(n19946) );
  OAI211_X1 U11831 ( .C1(n2954), .C2(n26614), .A(n19945), .B(n19946), .ZN(
        n19939) );
  OAI22_X1 U11836 ( .A1(n2952), .A2(n25678), .B1(n25676), .B2(n24635), .ZN(
        n19937) );
  OAI22_X1 U10530 ( .A1(n18363), .A2(n24588), .B1(n18332), .B2(n24652), .ZN(
        n18598) );
  OAI22_X1 U10531 ( .A1(n2196), .A2(net716477), .B1(net767232), .B2(n24651), 
        .ZN(n18597) );
  OAI22_X1 U10529 ( .A1(n2193), .A2(n18361), .B1(n2192), .B2(n18362), .ZN(
        n18599) );
  OAI22_X1 U10543 ( .A1(n2211), .A2(n18393), .B1(n2208), .B2(n18394), .ZN(
        n18616) );
  AOI21_X1 U10542 ( .B1(net767239), .B2(n17974), .A(n18616), .ZN(n18611) );
  OAI22_X1 U10541 ( .A1(n2205), .A2(n18390), .B1(n2190), .B2(n18318), .ZN(
        n18613) );
  OAI22_X1 U10540 ( .A1(n2209), .A2(n18387), .B1(n18388), .B2(n24649), .ZN(
        n18614) );
  AOI211_X1 U10539 ( .C1(net716405), .C2(n17984), .A(n18613), .B(n18614), .ZN(
        n18612) );
  OAI211_X1 U10538 ( .C1(n2212), .C2(n18382), .A(n18611), .B(n18612), .ZN(
        n18610) );
  AOI22_X1 U10545 ( .A1(net716417), .A2(n17975), .B1(net767235), .B2(n17985), 
        .ZN(n18617) );
  OAI21_X1 U10544 ( .B1(n2214), .B2(n18395), .A(n18617), .ZN(n18609) );
  OAI22_X1 U10547 ( .A1(n2206), .A2(n18400), .B1(n2189), .B2(n18401), .ZN(
        n18618) );
  OAI22_X1 U10532 ( .A1(n2195), .A2(n18369), .B1(net767237), .B2(n24650), .ZN(
        n18596) );
  OAI22_X1 U10389 ( .A1(n18363), .A2(n24589), .B1(n18332), .B2(n24662), .ZN(
        n18412) );
  OAI22_X1 U10390 ( .A1(n2052), .A2(net716477), .B1(net767232), .B2(n24661), 
        .ZN(n18411) );
  OAI22_X1 U10388 ( .A1(n2049), .A2(n18361), .B1(n2048), .B2(n18362), .ZN(
        n18413) );
  OAI22_X1 U10402 ( .A1(n2067), .A2(n18393), .B1(n2064), .B2(n18394), .ZN(
        n18431) );
  AOI21_X1 U10401 ( .B1(net767239), .B2(n17910), .A(n18431), .ZN(n18426) );
  OAI22_X1 U10400 ( .A1(n2061), .A2(n18390), .B1(n2046), .B2(n18318), .ZN(
        n18428) );
  OAI22_X1 U10399 ( .A1(n2065), .A2(n18387), .B1(n18388), .B2(n24659), .ZN(
        n18429) );
  AOI211_X1 U10398 ( .C1(net716405), .C2(n17920), .A(n18428), .B(n18429), .ZN(
        n18427) );
  OAI211_X1 U10397 ( .C1(n2068), .C2(n18382), .A(n18426), .B(n18427), .ZN(
        n18425) );
  AOI22_X1 U10404 ( .A1(net716417), .A2(n17911), .B1(net767235), .B2(n17921), 
        .ZN(n18432) );
  OAI21_X1 U10403 ( .B1(n2070), .B2(n18395), .A(n18432), .ZN(n18424) );
  OAI22_X1 U10406 ( .A1(n2062), .A2(n18400), .B1(n2045), .B2(n18401), .ZN(
        n18433) );
  OAI22_X1 U10391 ( .A1(n2051), .A2(n18369), .B1(net767237), .B2(n24660), .ZN(
        n18410) );
  OAI22_X1 U11084 ( .A1(n3108), .A2(n18346), .B1(n3107), .B2(net767172), .ZN(
        n19251) );
  OAI22_X1 U11079 ( .A1(n3089), .A2(n18401), .B1(net767232), .B2(n24627), .ZN(
        n19252) );
  OAI22_X1 U11075 ( .A1(n3103), .A2(net716477), .B1(net767237), .B2(n24628), 
        .ZN(n19253) );
  OAI22_X1 U11072 ( .A1(n3102), .A2(n18369), .B1(n3098), .B2(n18361), .ZN(
        n19254) );
  NOR4_X1 U11071 ( .A1(n19251), .A2(n19252), .A3(n19253), .A4(n19254), .ZN(
        n19232) );
  AOI22_X1 U11067 ( .A1(n18300), .A2(n24697), .B1(net767235), .B2(n18034), 
        .ZN(n19233) );
  NOR2_X1 U11060 ( .A1(n3124), .A2(n18394), .ZN(n19236) );
  OAI22_X1 U11057 ( .A1(n3131), .A2(n18382), .B1(n3130), .B2(n18393), .ZN(
        n19237) );
  AOI211_X1 U11056 ( .C1(n18022), .C2(net767239), .A(n19236), .B(n19237), .ZN(
        n19235) );
  AOI22_X1 U11063 ( .A1(n18307), .A2(n18035), .B1(net716405), .B2(n18033), 
        .ZN(n19234) );
  AOI22_X1 U11092 ( .A1(net767167), .A2(n24696), .B1(n18326), .B2(n18023), 
        .ZN(n19269) );
  AOI22_X1 U11097 ( .A1(net767238), .A2(n18021), .B1(net767171), .B2(n18027), 
        .ZN(n19268) );
  AOI22_X1 U11102 ( .A1(net716423), .A2(n18025), .B1(net767214), .B2(n18028), 
        .ZN(n19267) );
  AOI22_X1 U11111 ( .A1(n18372), .A2(n18032), .B1(n18373), .B2(n18031), .ZN(
        n19275) );
  AOI22_X1 U11105 ( .A1(n18330), .A2(n24695), .B1(n18331), .B2(n18026), .ZN(
        n19266) );
  OAI22_X1 U11417 ( .A1(n551), .A2(n19323), .B1(n550), .B2(n19324), .ZN(n19593) );
  AOI22_X1 U11416 ( .A1(n19327), .A2(n534), .B1(n19328), .B2(n536), .ZN(n19595) );
  NAND2_X1 U11415 ( .A1(n19530), .A2(n528), .ZN(n19596) );
  OAI211_X1 U11414 ( .C1(n543), .C2(n26785), .A(n19595), .B(n19596), .ZN(
        n19594) );
  AOI211_X1 U11413 ( .C1(n19320), .C2(n537), .A(n19593), .B(n19594), .ZN(
        n19587) );
  AOI22_X1 U11412 ( .A1(n25679), .A2(n529), .B1(n25666), .B2(n535), .ZN(n19588) );
  NOR2_X1 U11410 ( .A1(n549), .A2(n25677), .ZN(n19591) );
  OAI22_X1 U11409 ( .A1(n548), .A2(n25675), .B1(n25678), .B2(n24648), .ZN(
        n19592) );
  AOI211_X1 U11408 ( .C1(n524), .C2(n19348), .A(n19591), .B(n19592), .ZN(
        n19590) );
  AOI22_X1 U11411 ( .A1(n19344), .A2(n533), .B1(n19345), .B2(n530), .ZN(n19589) );
  AOI22_X1 U11428 ( .A1(n19336), .A2(n531), .B1(n19337), .B2(n17709), .ZN(
        n19601) );
  AOI22_X1 U11425 ( .A1(n24026), .A2(n526), .B1(n25682), .B2(n24762), .ZN(
        n19603) );
  AOI22_X1 U11423 ( .A1(n19308), .A2(n527), .B1(n23995), .B2(n24763), .ZN(
        n19597) );
  AOI22_X1 U11427 ( .A1(n24007), .A2(n17708), .B1(n25681), .B2(n17710), .ZN(
        n19602) );
  AOI22_X1 U11419 ( .A1(n19315), .A2(n17712), .B1(n25683), .B2(n17711), .ZN(
        n19600) );
  AOI22_X1 U11420 ( .A1(n23994), .A2(n24722), .B1(n19314), .B2(n538), .ZN(
        n19599) );
  AOI22_X1 U11422 ( .A1(n19318), .A2(n539), .B1(n19319), .B2(n525), .ZN(n19598) );
  OAI22_X1 U11998 ( .A1(n3108), .A2(n19350), .B1(n3107), .B2(n26614), .ZN(
        n20072) );
  OAI22_X1 U11993 ( .A1(n3089), .A2(n19396), .B1(n25677), .B2(n24627), .ZN(
        n20073) );
  OAI22_X1 U11989 ( .A1(n3103), .A2(n25678), .B1(n25675), .B2(n24628), .ZN(
        n20074) );
  OAI22_X1 U11986 ( .A1(n3102), .A2(n19370), .B1(n3098), .B2(n19365), .ZN(
        n20075) );
  NOR4_X1 U11985 ( .A1(n20072), .A2(n20073), .A3(n20074), .A4(n20075), .ZN(
        n20054) );
  AOI22_X1 U11980 ( .A1(n19308), .A2(n24697), .B1(n23995), .B2(n18034), .ZN(
        n20055) );
  NOR2_X1 U11973 ( .A1(n3124), .A2(n19389), .ZN(n20058) );
  OAI22_X1 U11970 ( .A1(n3131), .A2(n19378), .B1(n3130), .B2(n19388), .ZN(
        n20059) );
  AOI211_X1 U11969 ( .C1(n23994), .C2(n18022), .A(n20058), .B(n20059), .ZN(
        n20057) );
  AOI22_X1 U11976 ( .A1(n19315), .A2(n18035), .B1(n25683), .B2(n18033), .ZN(
        n20056) );
  AOI22_X1 U12020 ( .A1(n19336), .A2(n24695), .B1(n19337), .B2(n18026), .ZN(
        n20085) );
  AOI22_X1 U12027 ( .A1(n19372), .A2(n18032), .B1(n19373), .B2(n18031), .ZN(
        n20092) );
  AOI22_X1 U12006 ( .A1(n24026), .A2(n24696), .B1(n19333), .B2(n18023), .ZN(
        n20088) );
  AOI22_X1 U12012 ( .A1(n25674), .A2(n18021), .B1(n25680), .B2(n18027), .ZN(
        n20087) );
  AOI22_X1 U12017 ( .A1(n24007), .A2(n18025), .B1(n25681), .B2(n18028), .ZN(
        n20086) );
  OAI22_X1 U11669 ( .A1(n902), .A2(n19323), .B1(n901), .B2(n19324), .ZN(n19813) );
  AOI22_X1 U11668 ( .A1(n19327), .A2(n885), .B1(n19328), .B2(n887), .ZN(n19815) );
  NAND2_X1 U11667 ( .A1(n19530), .A2(n879), .ZN(n19816) );
  OAI211_X1 U11666 ( .C1(n894), .C2(n26785), .A(n19815), .B(n19816), .ZN(
        n19814) );
  AOI211_X1 U11665 ( .C1(n19320), .C2(n888), .A(n19813), .B(n19814), .ZN(
        n19807) );
  AOI22_X1 U11664 ( .A1(n25679), .A2(n880), .B1(n25667), .B2(n886), .ZN(n19808) );
  NOR2_X1 U11662 ( .A1(n900), .A2(n25677), .ZN(n19811) );
  OAI22_X1 U11661 ( .A1(n899), .A2(n25675), .B1(n25678), .B2(n24643), .ZN(
        n19812) );
  AOI211_X1 U11660 ( .C1(n875), .C2(n19348), .A(n19811), .B(n19812), .ZN(
        n19810) );
  AOI22_X1 U11663 ( .A1(n19344), .A2(n884), .B1(n19345), .B2(n881), .ZN(n19809) );
  AOI22_X1 U11680 ( .A1(n19336), .A2(n882), .B1(n19337), .B2(n17773), .ZN(
        n19821) );
  AOI22_X1 U11677 ( .A1(n24026), .A2(n877), .B1(n19333), .B2(n24752), .ZN(
        n19823) );
  AOI22_X1 U11675 ( .A1(n19308), .A2(n878), .B1(n23995), .B2(n24753), .ZN(
        n19817) );
  AOI22_X1 U11679 ( .A1(n24007), .A2(n17772), .B1(n19335), .B2(n17774), .ZN(
        n19822) );
  AOI22_X1 U11671 ( .A1(n19315), .A2(n17776), .B1(n25683), .B2(n17775), .ZN(
        n19820) );
  AOI22_X1 U11672 ( .A1(n23994), .A2(n24717), .B1(n19314), .B2(n889), .ZN(
        n19819) );
  AOI22_X1 U11674 ( .A1(n19318), .A2(n890), .B1(n19319), .B2(n876), .ZN(n19818) );
  OAI22_X1 U11719 ( .A1(n708), .A2(n19323), .B1(n707), .B2(n19324), .ZN(n19857) );
  AOI22_X1 U11718 ( .A1(n19327), .A2(n691), .B1(n19328), .B2(n693), .ZN(n19859) );
  NAND2_X1 U11717 ( .A1(n19530), .A2(n685), .ZN(n19860) );
  OAI211_X1 U11716 ( .C1(n700), .C2(n26785), .A(n19859), .B(n19860), .ZN(
        n19858) );
  AOI211_X1 U11715 ( .C1(n19320), .C2(n694), .A(n19857), .B(n19858), .ZN(
        n19851) );
  AOI22_X1 U11714 ( .A1(n25679), .A2(n686), .B1(n25667), .B2(n692), .ZN(n19852) );
  NOR2_X1 U11712 ( .A1(n706), .A2(n25677), .ZN(n19855) );
  OAI22_X1 U11711 ( .A1(n705), .A2(n25675), .B1(n25678), .B2(n24642), .ZN(
        n19856) );
  AOI211_X1 U11710 ( .C1(n681), .C2(n19348), .A(n19855), .B(n19856), .ZN(
        n19854) );
  AOI22_X1 U11713 ( .A1(n19344), .A2(n690), .B1(n19345), .B2(n687), .ZN(n19853) );
  AOI22_X1 U11730 ( .A1(n19336), .A2(n688), .B1(n19337), .B2(n17738), .ZN(
        n19865) );
  AOI22_X1 U11727 ( .A1(n24026), .A2(n683), .B1(n19333), .B2(n24750), .ZN(
        n19867) );
  AOI22_X1 U11725 ( .A1(n19308), .A2(n684), .B1(n23995), .B2(n24751), .ZN(
        n19861) );
  AOI22_X1 U11729 ( .A1(n24007), .A2(n17737), .B1(n19335), .B2(n17739), .ZN(
        n19866) );
  AOI22_X1 U11721 ( .A1(n19315), .A2(n17741), .B1(n25683), .B2(n17740), .ZN(
        n19864) );
  AOI22_X1 U11722 ( .A1(n23994), .A2(n24716), .B1(n19314), .B2(n695), .ZN(
        n19863) );
  AOI22_X1 U11724 ( .A1(n19318), .A2(n696), .B1(n19319), .B2(n682), .ZN(n19862) );
  OAI22_X1 U11018 ( .A1(n3063), .A2(n18346), .B1(n3062), .B2(net767172), .ZN(
        n19180) );
  OAI22_X1 U11017 ( .A1(n3053), .A2(n18401), .B1(n18367), .B2(n24631), .ZN(
        n19181) );
  OAI22_X1 U11016 ( .A1(n3060), .A2(net716477), .B1(net767237), .B2(n24632), 
        .ZN(n19182) );
  OAI22_X1 U11015 ( .A1(n3059), .A2(n18369), .B1(n3057), .B2(n18361), .ZN(
        n19183) );
  NOR4_X1 U11014 ( .A1(n19180), .A2(n19181), .A3(n19182), .A4(n19183), .ZN(
        n19173) );
  AOI22_X1 U11013 ( .A1(n18300), .A2(n24703), .B1(net767235), .B2(n17890), 
        .ZN(n19174) );
  NOR2_X1 U11011 ( .A1(n3072), .A2(n18394), .ZN(n19177) );
  OAI22_X1 U11010 ( .A1(n3076), .A2(n18382), .B1(n3075), .B2(n18393), .ZN(
        n19178) );
  AOI211_X1 U11009 ( .C1(n17878), .C2(net767239), .A(n19177), .B(n19178), .ZN(
        n19176) );
  AOI22_X1 U11012 ( .A1(n18307), .A2(n17891), .B1(net716405), .B2(n17889), 
        .ZN(n19175) );
  AOI22_X1 U11020 ( .A1(net767167), .A2(n24702), .B1(net716417), .B2(n17879), 
        .ZN(n19189) );
  AOI22_X1 U11021 ( .A1(net767238), .A2(n17877), .B1(net767171), .B2(n17883), 
        .ZN(n19188) );
  AOI22_X1 U11022 ( .A1(net716423), .A2(n17881), .B1(net767214), .B2(n17884), 
        .ZN(n19187) );
  AOI22_X1 U11025 ( .A1(n18372), .A2(n17888), .B1(n18373), .B2(n17887), .ZN(
        n19193) );
  AOI22_X1 U11023 ( .A1(n18330), .A2(n24701), .B1(n18331), .B2(n17882), .ZN(
        n19186) );
  OAI22_X1 U11442 ( .A1(n590), .A2(n19323), .B1(n589), .B2(n19324), .ZN(n19615) );
  AOI22_X1 U11441 ( .A1(n19327), .A2(n573), .B1(n19328), .B2(n575), .ZN(n19617) );
  NAND2_X1 U11440 ( .A1(n19530), .A2(n567), .ZN(n19618) );
  OAI211_X1 U11439 ( .C1(n582), .C2(n26785), .A(n19617), .B(n19618), .ZN(
        n19616) );
  AOI211_X1 U11438 ( .C1(n19320), .C2(n576), .A(n19615), .B(n19616), .ZN(
        n19609) );
  AOI22_X1 U11437 ( .A1(n25679), .A2(n568), .B1(n19351), .B2(n574), .ZN(n19610) );
  NOR2_X1 U11435 ( .A1(n588), .A2(n25677), .ZN(n19613) );
  OAI22_X1 U11434 ( .A1(n587), .A2(n25675), .B1(n25678), .B2(n24647), .ZN(
        n19614) );
  AOI211_X1 U11433 ( .C1(n563), .C2(n19348), .A(n19613), .B(n19614), .ZN(
        n19612) );
  AOI22_X1 U11436 ( .A1(n19344), .A2(n572), .B1(n19345), .B2(n569), .ZN(n19611) );
  AOI22_X1 U11453 ( .A1(n19336), .A2(n570), .B1(n19337), .B2(n17716), .ZN(
        n19623) );
  AOI22_X1 U11450 ( .A1(n24026), .A2(n565), .B1(n25682), .B2(n24760), .ZN(
        n19625) );
  AOI22_X1 U11448 ( .A1(n19308), .A2(n566), .B1(n23995), .B2(n24761), .ZN(
        n19619) );
  AOI22_X1 U11452 ( .A1(n24007), .A2(n17715), .B1(n19335), .B2(n17717), .ZN(
        n19624) );
  AOI22_X1 U11444 ( .A1(n19315), .A2(n17719), .B1(n25683), .B2(n17718), .ZN(
        n19622) );
  AOI22_X1 U11445 ( .A1(n23994), .A2(n24721), .B1(n19314), .B2(n577), .ZN(
        n19621) );
  AOI22_X1 U11447 ( .A1(n19318), .A2(n578), .B1(n19319), .B2(n564), .ZN(n19620) );
  OAI22_X1 U10996 ( .A1(n3027), .A2(n18346), .B1(n3026), .B2(net767172), .ZN(
        n19152) );
  OAI22_X1 U10995 ( .A1(n3017), .A2(n18401), .B1(net767232), .B2(n24633), .ZN(
        n19153) );
  OAI22_X1 U10994 ( .A1(n3024), .A2(net716477), .B1(net767237), .B2(n24634), 
        .ZN(n19154) );
  OAI22_X1 U10993 ( .A1(n3023), .A2(n18369), .B1(n3021), .B2(n18361), .ZN(
        n19155) );
  NOR4_X1 U10992 ( .A1(n19152), .A2(n19153), .A3(n19154), .A4(n19155), .ZN(
        n19145) );
  AOI22_X1 U10991 ( .A1(n18300), .A2(n24706), .B1(net767235), .B2(n17873), 
        .ZN(n19146) );
  NOR2_X1 U10989 ( .A1(n3036), .A2(n18394), .ZN(n19149) );
  OAI22_X1 U10988 ( .A1(n3040), .A2(n18382), .B1(n3039), .B2(n18393), .ZN(
        n19150) );
  AOI211_X1 U10987 ( .C1(n17861), .C2(net767239), .A(n19149), .B(n19150), .ZN(
        n19148) );
  AOI22_X1 U10990 ( .A1(n18307), .A2(n17874), .B1(net716405), .B2(n17872), 
        .ZN(n19147) );
  AOI22_X1 U10998 ( .A1(net767167), .A2(n24705), .B1(n18326), .B2(n17862), 
        .ZN(n19161) );
  AOI22_X1 U10999 ( .A1(net767238), .A2(n17860), .B1(net767171), .B2(n17866), 
        .ZN(n19160) );
  AOI22_X1 U11000 ( .A1(net716423), .A2(n17864), .B1(net767214), .B2(n17867), 
        .ZN(n19159) );
  AOI22_X1 U11003 ( .A1(n18372), .A2(n17871), .B1(n18373), .B2(n17870), .ZN(
        n19165) );
  AOI22_X1 U11001 ( .A1(n18330), .A2(n24704), .B1(n18331), .B2(n17865), .ZN(
        n19158) );
  AOI22_X1 U10933 ( .A1(n18372), .A2(n17837), .B1(n18373), .B2(n17836), .ZN(
        n19082) );
  AOI22_X1 U10931 ( .A1(n18330), .A2(n24709), .B1(n18331), .B2(n17831), .ZN(
        n19075) );
  OAI22_X1 U10515 ( .A1(n511), .A2(n18315), .B1(n510), .B2(n18316), .ZN(n18574) );
  AOI22_X1 U10514 ( .A1(net767173), .A2(n494), .B1(n18321), .B2(n496), .ZN(
        n18576) );
  NAND2_X1 U10513 ( .A1(n18529), .A2(n488), .ZN(n18577) );
  OAI211_X1 U10512 ( .C1(n503), .C2(net518461), .A(n18576), .B(n18577), .ZN(
        n18575) );
  AOI211_X1 U10511 ( .C1(n18312), .C2(n497), .A(n18574), .B(n18575), .ZN(
        n18567) );
  AOI22_X1 U10517 ( .A1(n18307), .A2(n17705), .B1(net716405), .B2(n17704), 
        .ZN(n18581) );
  AOI22_X1 U10518 ( .A1(net767239), .A2(n24723), .B1(n18306), .B2(n498), .ZN(
        n18580) );
  AOI22_X1 U10519 ( .A1(n18310), .A2(n499), .B1(n18311), .B2(n485), .ZN(n18579) );
  AOI22_X1 U10510 ( .A1(net716461), .A2(n489), .B1(n18347), .B2(n495), .ZN(
        n18568) );
  NOR2_X1 U10508 ( .A1(n509), .A2(net767232), .ZN(n18571) );
  OAI22_X1 U10507 ( .A1(n508), .A2(net767237), .B1(net716477), .B2(n24653), 
        .ZN(n18572) );
  AOI211_X1 U10506 ( .C1(n484), .C2(n18343), .A(n18571), .B(n18572), .ZN(
        n18570) );
  AOI22_X1 U10509 ( .A1(n18338), .A2(n493), .B1(n18339), .B2(n490), .ZN(n18569) );
  AOI22_X1 U10523 ( .A1(n18330), .A2(n491), .B1(n18331), .B2(n17702), .ZN(
        n18584) );
  AOI22_X1 U10521 ( .A1(net767167), .A2(n486), .B1(net716417), .B2(n24764), 
        .ZN(n18586) );
  AOI22_X1 U10520 ( .A1(n18300), .A2(n487), .B1(net767235), .B2(n24765), .ZN(
        n18578) );
  AOI22_X1 U10522 ( .A1(n18328), .A2(n17701), .B1(net767214), .B2(n17703), 
        .ZN(n18585) );
  AOI22_X1 U11190 ( .A1(n25682), .A2(n17896), .B1(n23995), .B2(n17906), .ZN(
        n19391) );
  OAI21_X1 U11189 ( .B1(n2034), .B2(n19390), .A(n19391), .ZN(n19376) );
  OAI22_X1 U11188 ( .A1(n2031), .A2(n19388), .B1(n2028), .B2(n19389), .ZN(
        n19387) );
  AOI21_X1 U11187 ( .B1(n23994), .B2(n17895), .A(n19387), .ZN(n19379) );
  OAI22_X1 U11186 ( .A1(n2025), .A2(n19385), .B1(n2010), .B2(n19326), .ZN(
        n19381) );
  OAI22_X1 U11185 ( .A1(n2029), .A2(n19383), .B1(n19384), .B2(n24663), .ZN(
        n19382) );
  AOI211_X1 U11184 ( .C1(n25683), .C2(n17905), .A(n19381), .B(n19382), .ZN(
        n19380) );
  OAI211_X1 U11183 ( .C1(n2032), .C2(n19378), .A(n19379), .B(n19380), .ZN(
        n19377) );
  AOI211_X1 U11182 ( .C1(n24026), .C2(n24724), .A(n19376), .B(n19377), .ZN(
        n19375) );
  OAI22_X1 U11193 ( .A1(n2026), .A2(n19395), .B1(n2009), .B2(n19396), .ZN(
        n19394) );
  AOI21_X1 U11192 ( .B1(n25674), .B2(n17894), .A(n19394), .ZN(n19374) );
  OAI22_X1 U11175 ( .A1(n2015), .A2(n19370), .B1(n25676), .B2(n24664), .ZN(
        n19361) );
  OAI22_X1 U11174 ( .A1(n2016), .A2(n25678), .B1(n25677), .B2(n24665), .ZN(
        n19362) );
  OAI22_X1 U11173 ( .A1(n19367), .A2(n24590), .B1(n19338), .B2(n24666), .ZN(
        n19363) );
  OAI22_X1 U11172 ( .A1(n2013), .A2(n19365), .B1(n2012), .B2(n19366), .ZN(
        n19364) );
  NOR4_X1 U11171 ( .A1(n19361), .A2(n19362), .A3(n19363), .A4(n19364), .ZN(
        n19360) );
  AOI22_X1 U11180 ( .A1(n19334), .A2(n17897), .B1(n25681), .B2(n17900), .ZN(
        n19357) );
  AOI22_X1 U11177 ( .A1(n25679), .A2(n24598), .B1(n25667), .B2(n24790), .ZN(
        n19358) );
  AOI22_X1 U11176 ( .A1(n19372), .A2(n17904), .B1(n19373), .B2(n17903), .ZN(
        n19359) );
  NOR2_X1 U11292 ( .A1(n2154), .A2(n19326), .ZN(n19489) );
  OAI22_X1 U11291 ( .A1(n2169), .A2(n19385), .B1(n2170), .B2(n19395), .ZN(
        n19490) );
  AOI22_X1 U11288 ( .A1(n25674), .A2(n17958), .B1(n19332), .B2(n24727), .ZN(
        n19482) );
  AOI22_X1 U11286 ( .A1(n25682), .A2(n17960), .B1(n19308), .B2(n24728), .ZN(
        n19483) );
  AOI22_X1 U11284 ( .A1(n23995), .A2(n17969), .B1(n19318), .B2(n24804), .ZN(
        n19484) );
  AOI22_X1 U11282 ( .A1(n19319), .A2(n24793), .B1(n23994), .B2(n17959), .ZN(
        n19485) );
  NAND4_X1 U11281 ( .A1(n19482), .A2(n19483), .A3(n19484), .A4(n19485), .ZN(
        n19473) );
  OAI22_X1 U11280 ( .A1(n2153), .A2(n19396), .B1(n2173), .B2(n19383), .ZN(
        n19474) );
  OAI22_X1 U11279 ( .A1(n2172), .A2(n19389), .B1(n24615), .B2(n24777), .ZN(
        n19475) );
  AOI22_X1 U11278 ( .A1(n19315), .A2(n17970), .B1(n19372), .B2(n17967), .ZN(
        n19478) );
  NAND2_X1 U11277 ( .A1(n19373), .A2(n17966), .ZN(n19479) );
  OAI211_X1 U11276 ( .C1(n2162), .C2(n26614), .A(n19478), .B(n19479), .ZN(
        n19476) );
  NOR4_X1 U11275 ( .A1(n19473), .A2(n19474), .A3(n19475), .A4(n19476), .ZN(
        n19472) );
  AOI22_X1 U11296 ( .A1(n19334), .A2(n17961), .B1(n19337), .B2(n17962), .ZN(
        n19493) );
  AOI22_X1 U11293 ( .A1(n25681), .A2(n17963), .B1(n25680), .B2(n14393), .ZN(
        n19470) );
  AOI22_X1 U11294 ( .A1(n24619), .A2(n17965), .B1(n24591), .B2(n17964), .ZN(
        n19469) );
  AOI22_X1 U11376 ( .A1(n25682), .A2(n17975), .B1(n23995), .B2(n17985), .ZN(
        n19558) );
  OAI21_X1 U11375 ( .B1(n2214), .B2(n19390), .A(n19558), .ZN(n19551) );
  OAI22_X1 U11374 ( .A1(n2211), .A2(n19388), .B1(n2208), .B2(n19389), .ZN(
        n19557) );
  AOI21_X1 U11373 ( .B1(n23994), .B2(n17974), .A(n19557), .ZN(n19553) );
  OAI22_X1 U11372 ( .A1(n2205), .A2(n19385), .B1(n2190), .B2(n19326), .ZN(
        n19555) );
  OAI22_X1 U11371 ( .A1(n2209), .A2(n19383), .B1(n19384), .B2(n24649), .ZN(
        n19556) );
  AOI211_X1 U11370 ( .C1(n25683), .C2(n17984), .A(n19555), .B(n19556), .ZN(
        n19554) );
  OAI211_X1 U11369 ( .C1(n2212), .C2(n19378), .A(n19553), .B(n19554), .ZN(
        n19552) );
  AOI211_X1 U11368 ( .C1(n24026), .C2(n24725), .A(n19551), .B(n19552), .ZN(
        n19550) );
  OAI22_X1 U11379 ( .A1(n2206), .A2(n19395), .B1(n2189), .B2(n19396), .ZN(
        n19559) );
  AOI21_X1 U11378 ( .B1(n25674), .B2(n17973), .A(n19559), .ZN(n19549) );
  OAI22_X1 U11361 ( .A1(n2195), .A2(n19370), .B1(n25675), .B2(n24650), .ZN(
        n19545) );
  OAI22_X1 U11360 ( .A1(n2196), .A2(n25678), .B1(n25677), .B2(n24651), .ZN(
        n19546) );
  OAI22_X1 U11359 ( .A1(n19367), .A2(n24588), .B1(n19338), .B2(n24652), .ZN(
        n19547) );
  OAI22_X1 U11358 ( .A1(n2193), .A2(n19365), .B1(n2192), .B2(n19366), .ZN(
        n19548) );
  NOR4_X1 U11357 ( .A1(n19545), .A2(n19546), .A3(n19547), .A4(n19548), .ZN(
        n19544) );
  AOI22_X1 U11366 ( .A1(n19334), .A2(n17976), .B1(n25681), .B2(n17979), .ZN(
        n19541) );
  AOI22_X1 U11363 ( .A1(n25679), .A2(n24599), .B1(n25666), .B2(n24791), .ZN(
        n19542) );
  AOI22_X1 U11362 ( .A1(n19372), .A2(n17983), .B1(n19373), .B2(n17982), .ZN(
        n19543) );
  AOI22_X1 U11216 ( .A1(n25682), .A2(n17911), .B1(n23995), .B2(n17921), .ZN(
        n19417) );
  OAI21_X1 U11215 ( .B1(n2070), .B2(n19390), .A(n19417), .ZN(n19410) );
  OAI22_X1 U11214 ( .A1(n2067), .A2(n19388), .B1(n2064), .B2(n19389), .ZN(
        n19416) );
  AOI21_X1 U11213 ( .B1(n23994), .B2(n17910), .A(n19416), .ZN(n19412) );
  OAI22_X1 U11212 ( .A1(n2061), .A2(n19385), .B1(n2046), .B2(n19326), .ZN(
        n19414) );
  OAI22_X1 U11211 ( .A1(n2065), .A2(n19383), .B1(n19384), .B2(n24659), .ZN(
        n19415) );
  AOI211_X1 U11210 ( .C1(n25683), .C2(n17920), .A(n19414), .B(n19415), .ZN(
        n19413) );
  OAI211_X1 U11209 ( .C1(n2068), .C2(n19378), .A(n19412), .B(n19413), .ZN(
        n19411) );
  AOI211_X1 U11208 ( .C1(n24026), .C2(n24726), .A(n19410), .B(n19411), .ZN(
        n19409) );
  OAI22_X1 U11219 ( .A1(n2062), .A2(n19395), .B1(n2045), .B2(n19396), .ZN(
        n19418) );
  AOI21_X1 U11218 ( .B1(n25674), .B2(n17909), .A(n19418), .ZN(n19408) );
  OAI22_X1 U11201 ( .A1(n2051), .A2(n19370), .B1(n25675), .B2(n24660), .ZN(
        n19404) );
  OAI22_X1 U11200 ( .A1(n2052), .A2(n25678), .B1(n25677), .B2(n24661), .ZN(
        n19405) );
  OAI22_X1 U11199 ( .A1(n19367), .A2(n24589), .B1(n19338), .B2(n24662), .ZN(
        n19406) );
  OAI22_X1 U11198 ( .A1(n2049), .A2(n19365), .B1(n2048), .B2(n19366), .ZN(
        n19407) );
  NOR4_X1 U11197 ( .A1(n19404), .A2(n19405), .A3(n19406), .A4(n19407), .ZN(
        n19403) );
  AOI22_X1 U11206 ( .A1(n19334), .A2(n17912), .B1(n25681), .B2(n17915), .ZN(
        n19400) );
  AOI22_X1 U11203 ( .A1(n25679), .A2(n24600), .B1(n25667), .B2(n24792), .ZN(
        n19401) );
  AOI22_X1 U11202 ( .A1(n19372), .A2(n17919), .B1(n19373), .B2(n17918), .ZN(
        n19402) );
  OAI22_X1 U11860 ( .A1(n2991), .A2(n19350), .B1(n2990), .B2(n26614), .ZN(
        n19964) );
  OAI22_X1 U11859 ( .A1(n2981), .A2(n19396), .B1(n25677), .B2(n24620), .ZN(
        n19965) );
  OAI22_X1 U11858 ( .A1(n2988), .A2(n25678), .B1(n25676), .B2(n24621), .ZN(
        n19966) );
  OAI22_X1 U11857 ( .A1(n2987), .A2(n19370), .B1(n2985), .B2(n19365), .ZN(
        n19967) );
  NOR4_X1 U11856 ( .A1(n19964), .A2(n19965), .A3(n19966), .A4(n19967), .ZN(
        n19958) );
  AOI22_X1 U11854 ( .A1(n19308), .A2(n24684), .B1(n23995), .B2(n17856), .ZN(
        n19959) );
  AOI22_X1 U11853 ( .A1(n19315), .A2(n17857), .B1(n25683), .B2(n17855), .ZN(
        n19960) );
  NOR2_X1 U11852 ( .A1(n3000), .A2(n19389), .ZN(n19962) );
  OAI22_X1 U11851 ( .A1(n3004), .A2(n19378), .B1(n3003), .B2(n19388), .ZN(
        n19963) );
  AOI211_X1 U11850 ( .C1(n23994), .C2(n17844), .A(n19962), .B(n19963), .ZN(
        n19961) );
  AOI22_X1 U11864 ( .A1(n25674), .A2(n17843), .B1(n25680), .B2(n17849), .ZN(
        n19970) );
  AOI22_X1 U11862 ( .A1(n19332), .A2(n24683), .B1(n25682), .B2(n17845), .ZN(
        n19971) );
  AOI22_X1 U11865 ( .A1(n24007), .A2(n17847), .B1(n19335), .B2(n17850), .ZN(
        n19969) );
  OAI22_X1 U10630 ( .A1(n629), .A2(n18315), .B1(n628), .B2(n18316), .ZN(n18713) );
  AOI22_X1 U10629 ( .A1(net767173), .A2(n612), .B1(n18321), .B2(n614), .ZN(
        n18715) );
  NAND2_X1 U10628 ( .A1(n18529), .A2(n606), .ZN(n18716) );
  OAI211_X1 U10627 ( .C1(n621), .C2(net518461), .A(n18715), .B(n18716), .ZN(
        n18714) );
  AOI211_X1 U10626 ( .C1(n18312), .C2(n615), .A(n18713), .B(n18714), .ZN(
        n18706) );
  AOI22_X1 U10632 ( .A1(n18307), .A2(n17727), .B1(net716405), .B2(n17726), 
        .ZN(n18720) );
  AOI22_X1 U10633 ( .A1(net767239), .A2(n24693), .B1(n18306), .B2(n616), .ZN(
        n18719) );
  AOI22_X1 U10634 ( .A1(n18310), .A2(n617), .B1(n18311), .B2(n603), .ZN(n18718) );
  AOI22_X1 U10625 ( .A1(net716461), .A2(n607), .B1(n18347), .B2(n613), .ZN(
        n18707) );
  NOR2_X1 U10623 ( .A1(n627), .A2(net767232), .ZN(n18710) );
  OAI22_X1 U10622 ( .A1(n626), .A2(net767237), .B1(net716477), .B2(n24625), 
        .ZN(n18711) );
  AOI211_X1 U10621 ( .C1(n602), .C2(n18343), .A(n18710), .B(n18711), .ZN(
        n18709) );
  AOI22_X1 U10624 ( .A1(n18338), .A2(n611), .B1(n18339), .B2(n608), .ZN(n18708) );
  AOI22_X1 U10638 ( .A1(n18330), .A2(n609), .B1(n18331), .B2(n17724), .ZN(
        n18723) );
  AOI22_X1 U10636 ( .A1(n18325), .A2(n604), .B1(net716417), .B2(n24743), .ZN(
        n18725) );
  AOI22_X1 U10635 ( .A1(n18300), .A2(n605), .B1(net767235), .B2(n24744), .ZN(
        n18717) );
  AOI22_X1 U10637 ( .A1(net716423), .A2(n17723), .B1(net767214), .B2(n17725), 
        .ZN(n18724) );
  OAI22_X1 U11805 ( .A1(n2919), .A2(n19350), .B1(n2918), .B2(n26614), .ZN(
        n19922) );
  OAI22_X1 U11804 ( .A1(n2909), .A2(n19396), .B1(n25677), .B2(n24637), .ZN(
        n19923) );
  OAI22_X1 U11803 ( .A1(n2916), .A2(n25678), .B1(n25675), .B2(n24638), .ZN(
        n19924) );
  OAI22_X1 U11802 ( .A1(n2915), .A2(n19370), .B1(n2913), .B2(n19365), .ZN(
        n19925) );
  NOR4_X1 U11801 ( .A1(n19922), .A2(n19923), .A3(n19924), .A4(n19925), .ZN(
        n19916) );
  AOI22_X1 U11807 ( .A1(n24026), .A2(n24710), .B1(n25682), .B2(n17828), .ZN(
        n19929) );
  AOI22_X1 U11809 ( .A1(n25674), .A2(n17826), .B1(n25680), .B2(n17832), .ZN(
        n19928) );
  AOI22_X1 U11810 ( .A1(n24007), .A2(n17830), .B1(n19335), .B2(n17833), .ZN(
        n19927) );
  AOI22_X1 U11799 ( .A1(n19308), .A2(n24711), .B1(n23995), .B2(n17839), .ZN(
        n19917) );
  NOR2_X1 U11797 ( .A1(n2928), .A2(n19389), .ZN(n19920) );
  OAI22_X1 U11796 ( .A1(n2932), .A2(n19378), .B1(n2931), .B2(n19388), .ZN(
        n19921) );
  AOI211_X1 U11795 ( .C1(n23994), .C2(n17827), .A(n19920), .B(n19921), .ZN(
        n19919) );
  AOI22_X1 U11798 ( .A1(n19315), .A2(n17840), .B1(n25683), .B2(n17838), .ZN(
        n19918) );
  AOI22_X1 U10946 ( .A1(n18300), .A2(n996), .B1(net767235), .B2(n17805), .ZN(
        n19094) );
  AOI22_X1 U10943 ( .A1(n18310), .A2(n24708), .B1(n18311), .B2(n994), .ZN(
        n19095) );
  AOI22_X1 U10941 ( .A1(net767239), .A2(n17794), .B1(n18306), .B2(n24747), 
        .ZN(n19096) );
  AOI22_X1 U10940 ( .A1(n18307), .A2(n17806), .B1(net716405), .B2(n17804), 
        .ZN(n19097) );
  NAND4_X1 U10939 ( .A1(n19094), .A2(n19095), .A3(n19096), .A4(n19097), .ZN(
        n19093) );
  AOI22_X1 U10949 ( .A1(n18343), .A2(n993), .B1(net716491), .B2(n17801), .ZN(
        n19100) );
  NAND2_X1 U10948 ( .A1(net716461), .A2(n998), .ZN(n19101) );
  OAI211_X1 U10947 ( .C1(n2954), .C2(net767172), .A(n19100), .B(n19101), .ZN(
        n19092) );
  OAI22_X1 U10951 ( .A1(n2951), .A2(n18369), .B1(n18361), .B2(n24636), .ZN(
        n19091) );
  AOI22_X1 U10954 ( .A1(net767167), .A2(n995), .B1(n18326), .B2(n17795), .ZN(
        n19107) );
  AOI22_X1 U10957 ( .A1(n18330), .A2(n24707), .B1(n18331), .B2(n14402), .ZN(
        n19104) );
  AOI22_X1 U10956 ( .A1(net716423), .A2(n17797), .B1(net767214), .B2(n17799), 
        .ZN(n19105) );
  AOI22_X1 U10955 ( .A1(net767238), .A2(n17793), .B1(net767171), .B2(n17798), 
        .ZN(n19106) );
  AOI22_X1 U10959 ( .A1(n18372), .A2(n17803), .B1(n18373), .B2(n17802), .ZN(
        n19110) );
  OAI22_X1 U10952 ( .A1(n2952), .A2(net716477), .B1(net767237), .B2(n24635), 
        .ZN(n19090) );
  OAI22_X1 U11749 ( .A1(n981), .A2(n19323), .B1(n980), .B2(n19324), .ZN(n19879) );
  AOI22_X1 U11745 ( .A1(n19327), .A2(n964), .B1(n19328), .B2(n966), .ZN(n19881) );
  NAND2_X1 U11744 ( .A1(n19530), .A2(n958), .ZN(n19882) );
  OAI211_X1 U11743 ( .C1(n973), .C2(n26785), .A(n19881), .B(n19882), .ZN(
        n19880) );
  AOI211_X1 U11742 ( .C1(n19320), .C2(n967), .A(n19879), .B(n19880), .ZN(
        n19873) );
  AOI22_X1 U11741 ( .A1(n25679), .A2(n959), .B1(n25667), .B2(n965), .ZN(n19874) );
  NOR2_X1 U11737 ( .A1(n979), .A2(n25677), .ZN(n19877) );
  OAI22_X1 U11736 ( .A1(n978), .A2(n25675), .B1(n25678), .B2(n24641), .ZN(
        n19878) );
  AOI211_X1 U11735 ( .C1(n954), .C2(n19348), .A(n19877), .B(n19878), .ZN(
        n19876) );
  AOI22_X1 U11738 ( .A1(n19344), .A2(n963), .B1(n19345), .B2(n960), .ZN(n19875) );
  AOI22_X1 U11763 ( .A1(n19336), .A2(n961), .B1(n19337), .B2(n17787), .ZN(
        n19887) );
  AOI22_X1 U11760 ( .A1(n24026), .A2(n956), .B1(n19333), .B2(n24748), .ZN(
        n19889) );
  AOI22_X1 U11758 ( .A1(n19308), .A2(n957), .B1(n23995), .B2(n24749), .ZN(
        n19883) );
  AOI22_X1 U11762 ( .A1(n24007), .A2(n17786), .B1(n19335), .B2(n17788), .ZN(
        n19888) );
  AOI22_X1 U11754 ( .A1(n19315), .A2(n17790), .B1(n25683), .B2(n17789), .ZN(
        n19886) );
  AOI22_X1 U11755 ( .A1(n23994), .A2(n24715), .B1(n19314), .B2(n968), .ZN(
        n19885) );
  AOI22_X1 U11757 ( .A1(n19318), .A2(n969), .B1(n19319), .B2(n955), .ZN(n19884) );
  OAI22_X1 U11467 ( .A1(n629), .A2(n19323), .B1(n628), .B2(n19324), .ZN(n19637) );
  AOI22_X1 U11466 ( .A1(n19327), .A2(n612), .B1(n19328), .B2(n614), .ZN(n19639) );
  NAND2_X1 U11465 ( .A1(n19530), .A2(n606), .ZN(n19640) );
  OAI211_X1 U11464 ( .C1(n621), .C2(n26785), .A(n19639), .B(n19640), .ZN(
        n19638) );
  AOI211_X1 U11463 ( .C1(n19320), .C2(n615), .A(n19637), .B(n19638), .ZN(
        n19631) );
  AOI22_X1 U11462 ( .A1(n25679), .A2(n607), .B1(n19351), .B2(n613), .ZN(n19632) );
  NOR2_X1 U11460 ( .A1(n627), .A2(n25677), .ZN(n19635) );
  OAI22_X1 U11459 ( .A1(n626), .A2(n25676), .B1(n25678), .B2(n24625), .ZN(
        n19636) );
  AOI211_X1 U11458 ( .C1(n602), .C2(n19348), .A(n19635), .B(n19636), .ZN(
        n19634) );
  AOI22_X1 U11461 ( .A1(n19344), .A2(n611), .B1(n19345), .B2(n608), .ZN(n19633) );
  AOI22_X1 U11478 ( .A1(n19336), .A2(n609), .B1(n19337), .B2(n17724), .ZN(
        n19645) );
  AOI22_X1 U11475 ( .A1(n24026), .A2(n604), .B1(n19333), .B2(n24743), .ZN(
        n19647) );
  AOI22_X1 U11473 ( .A1(n19308), .A2(n605), .B1(n23995), .B2(n24744), .ZN(
        n19641) );
  AOI22_X1 U11477 ( .A1(n24007), .A2(n17723), .B1(n25681), .B2(n17725), .ZN(
        n19646) );
  AOI22_X1 U11469 ( .A1(n19315), .A2(n17727), .B1(n25683), .B2(n17726), .ZN(
        n19644) );
  AOI22_X1 U11470 ( .A1(n23994), .A2(n24693), .B1(n19314), .B2(n616), .ZN(
        n19643) );
  AOI22_X1 U11472 ( .A1(n19318), .A2(n617), .B1(n19319), .B2(n603), .ZN(n19642) );
  NAND2_X1 U10139 ( .A1(n18131), .A2(n18135), .ZN(n18190) );
  OAI21_X1 U10138 ( .B1(net741565), .B2(net518455), .A(n18190), .ZN(
        \cu_inst/EX/DFF_10/N3 ) );
  NAND2_X1 U10137 ( .A1(net710387), .A2(n18190), .ZN(\cu_inst/EX/DFF_11/N3 )
         );
  AOI22_X1 U13796 ( .A1(n23997), .A2(n25616), .B1(n25082), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_16/N3 ) );
  AOI22_X1 U13643 ( .A1(n24024), .A2(n25618), .B1(n24861), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_17/N3 ) );
  AOI22_X1 U13593 ( .A1(n24022), .A2(n26768), .B1(n24876), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_16/N3 ) );
  AOI22_X1 U13749 ( .A1(n24014), .A2(n26773), .B1(n24852), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_10/N3 ) );
  AOI22_X1 U13626 ( .A1(n24024), .A2(n25634), .B1(n24867), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_25/N3 ) );
  AOI22_X1 U13574 ( .A1(n24022), .A2(n26758), .B1(n24883), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_25/N3 ) );
  AOI22_X1 U13738 ( .A1(n24014), .A2(n26768), .B1(n970), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_16/N3 ) );
  AOI22_X1 U13645 ( .A1(n24024), .A2(n25616), .B1(n24860), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_16/N3 ) );
  AOI22_X1 U13737 ( .A1(n24014), .A2(n26767), .B1(n697), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_17/N3 ) );
  AOI22_X1 U13654 ( .A1(n24024), .A2(n25604), .B1(n2719), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_1/N3 ) );
  AOI22_X1 U13721 ( .A1(n24014), .A2(n26753), .B1(n25036), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_3/N3 ) );
  AOI22_X1 U13653 ( .A1(n24024), .A2(n25606), .B1(n3079), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_10/N3 ) );
  AOI22_X1 U13688 ( .A1(n24013), .A2(n25617), .B1(n971), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_16/N3 ) );
  AOI22_X1 U13535 ( .A1(n24012), .A2(n25617), .B1(n972), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_16/N3 ) );
  AOI22_X1 U13777 ( .A1(n23997), .A2(n25634), .B1(n25089), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_25/N3 ) );
  AOI22_X1 U13601 ( .A1(n24022), .A2(n26773), .B1(n3078), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_10/N3 ) );
  AOI22_X1 U13804 ( .A1(n23997), .A2(n25606), .B1(n3075), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_10/N3 ) );
  AOI22_X1 U13518 ( .A1(n24012), .A2(n25645), .B1(n24889), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_3/N3 ) );
  AOI22_X1 U13671 ( .A1(n24013), .A2(n25645), .B1(n24844), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_3/N3 ) );
  AOI22_X1 U13591 ( .A1(n24022), .A2(n26767), .B1(n24877), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_17/N3 ) );
  AOI22_X1 U13544 ( .A1(n24012), .A2(n25609), .B1(n25101), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_11/N3 ) );
  AOI22_X1 U13546 ( .A1(n24012), .A2(n25607), .B1(n25100), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_10/N3 ) );
  AOI22_X1 U13699 ( .A1(n24013), .A2(n25607), .B1(n25273), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_10/N3 ) );
  AOI22_X1 U13805 ( .A1(n23997), .A2(n25604), .B1(n2715), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_1/N3 ) );
  AOI22_X1 U13516 ( .A1(n24012), .A2(n25649), .B1(n464), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_31/N3 ) );
  AOI22_X1 U13697 ( .A1(n24013), .A2(n25609), .B1(n25274), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_11/N3 ) );
  AOI22_X1 U13747 ( .A1(n24014), .A2(n26772), .B1(n24853), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_11/N3 ) );
  AOI22_X1 U13731 ( .A1(n24014), .A2(n26762), .B1(n735), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_21/N3 ) );
  AOI22_X1 U13727 ( .A1(n24014), .A2(n26758), .B1(n388), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_25/N3 ) );
  AOI22_X1 U13677 ( .A1(n24013), .A2(n25635), .B1(n389), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_25/N3 ) );
  AOI22_X1 U13524 ( .A1(n24012), .A2(n25635), .B1(n390), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_25/N3 ) );
  AOI22_X1 U13800 ( .A1(n23997), .A2(n25610), .B1(n25081), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_13/N3 ) );
  AOI22_X1 U13649 ( .A1(n24024), .A2(n25610), .B1(n24859), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_13/N3 ) );
  AOI22_X1 U13597 ( .A1(n24022), .A2(n26771), .B1(n24875), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_13/N3 ) );
  AOI22_X1 U13521 ( .A1(n24012), .A2(n25641), .B1(n542), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_28/N3 ) );
  AOI22_X1 U13674 ( .A1(n24013), .A2(n25641), .B1(n541), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_28/N3 ) );
  AOI22_X1 U13743 ( .A1(n24014), .A2(n26771), .B1(n24854), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_13/N3 ) );
  AOI22_X1 U13693 ( .A1(n24013), .A2(n25611), .B1(n24858), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_13/N3 ) );
  AOI22_X1 U13540 ( .A1(n24012), .A2(n25611), .B1(n25102), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_13/N3 ) );
  AOI22_X1 U13600 ( .A1(n24022), .A2(n26772), .B1(n3042), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_11/N3 ) );
  AOI22_X1 U13652 ( .A1(n24024), .A2(n25608), .B1(n3043), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_11/N3 ) );
  AOI22_X1 U13803 ( .A1(n23997), .A2(n25608), .B1(n3039), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_11/N3 ) );
  AOI22_X1 U13724 ( .A1(n24014), .A2(n26755), .B1(n540), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_28/N3 ) );
  AOI22_X1 U13580 ( .A1(n24022), .A2(n26761), .B1(net741196), .B2(n20613), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_14/DFF_22/N3 ) );
  AOI22_X1 U13632 ( .A1(n24024), .A2(net717153), .B1(net741214), .B2(n20632), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_13/DFF_22/N3 ) );
  AOI22_X1 U13526 ( .A1(n24012), .A2(n25631), .B1(n775), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_23/N3 ) );
  AOI22_X1 U13568 ( .A1(n24022), .A2(n26755), .B1(n24886), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_28/N3 ) );
  AOI22_X1 U13620 ( .A1(n24024), .A2(n25640), .B1(n24870), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_28/N3 ) );
  AOI22_X1 U13534 ( .A1(n24012), .A2(n25619), .B1(n699), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_17/N3 ) );
  AOI22_X1 U13798 ( .A1(n23997), .A2(n25614), .B1(n2895), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_15/N3 ) );
  AOI22_X1 U13647 ( .A1(n24024), .A2(n25614), .B1(n2899), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_15/N3 ) );
  AOI22_X1 U13595 ( .A1(n24022), .A2(n26769), .B1(n2898), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_15/N3 ) );
  AOI22_X1 U13771 ( .A1(n23997), .A2(n25640), .B1(n25092), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_28/N3 ) );
  AOI22_X1 U13789 ( .A1(n23997), .A2(n25624), .B1(n2319), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_2/N3 ) );
  AOI22_X1 U13638 ( .A1(n24024), .A2(n25624), .B1(n2323), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_2/N3 ) );
  AOI22_X1 U13739 ( .A1(n24014), .A2(n26769), .B1(n24856), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_15/N3 ) );
  AOI22_X1 U13689 ( .A1(n24013), .A2(n25615), .B1(n25276), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_15/N3 ) );
  AOI22_X1 U13536 ( .A1(n24012), .A2(n25615), .B1(n25104), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_15/N3 ) );
  AOI22_X1 U13586 ( .A1(n24022), .A2(n26764), .B1(n2322), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_2/N3 ) );
  AOI22_X1 U13764 ( .A1(n23997), .A2(n25648), .B1(n25095), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_31/N3 ) );
  AOI22_X1 U13613 ( .A1(n24024), .A2(n25648), .B1(n24873), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_31/N3 ) );
  AOI22_X1 U13561 ( .A1(n24022), .A2(n26751), .B1(n24655), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_31/N3 ) );
  AOI22_X1 U13530 ( .A1(n24012), .A2(n25625), .B1(n25306), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_2/N3 ) );
  AOI22_X1 U13683 ( .A1(n24013), .A2(n25625), .B1(n25313), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_2/N3 ) );
  AOI22_X1 U13719 ( .A1(n24014), .A2(n26751), .B1(n462), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_31/N3 ) );
  AOI22_X1 U13669 ( .A1(n24013), .A2(n25649), .B1(n463), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_31/N3 ) );
  AOI22_X1 U13733 ( .A1(n24014), .A2(n26764), .B1(n25284), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_2/N3 ) );
  AOI22_X1 U13783 ( .A1(n23997), .A2(net717153), .B1(net740970), .B2(n20686), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_10/DFF_22/N3 ) );
  AOI22_X1 U13602 ( .A1(n24022), .A2(n26774), .B1(n2718), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_1/N3 ) );
  AOI22_X1 U13715 ( .A1(n24014), .A2(n26749), .B1(n25097), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_5/N3 ) );
  AOI22_X1 U13678 ( .A1(n24013), .A2(n25633), .B1(n659), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_24/N3 ) );
  AOI22_X1 U13665 ( .A1(n24013), .A2(n25653), .B1(n25279), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_5/N3 ) );
  AOI22_X1 U13511 ( .A1(n24012), .A2(n25653), .B1(n25269), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_5/N3 ) );
  AOI22_X1 U13582 ( .A1(n24022), .A2(n26762), .B1(n24880), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_21/N3 ) );
  AOI22_X1 U13559 ( .A1(n24022), .A2(n26749), .B1(n2142), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_5/N3 ) );
  AOI22_X1 U13611 ( .A1(n24024), .A2(n25652), .B1(n2143), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_5/N3 ) );
  AOI22_X1 U13762 ( .A1(n23997), .A2(n25652), .B1(n2139), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_5/N3 ) );
  AOI22_X1 U13528 ( .A1(n24012), .A2(n25628), .B1(n737), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_21/N3 ) );
  AOI22_X1 U13681 ( .A1(n24013), .A2(n25628), .B1(n736), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_21/N3 ) );
  AOI22_X1 U13550 ( .A1(n24012), .A2(n25603), .B1(n25098), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_0/N3 ) );
  AOI22_X1 U13703 ( .A1(n24013), .A2(n25603), .B1(n25271), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_0/N3 ) );
  AOI22_X1 U13753 ( .A1(n24014), .A2(n26775), .B1(n24850), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_0/N3 ) );
  AOI22_X1 U13728 ( .A1(n24014), .A2(n26759), .B1(n658), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_24/N3 ) );
  AOI22_X1 U13525 ( .A1(n24012), .A2(n25633), .B1(n660), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_24/N3 ) );
  AOI22_X1 U13634 ( .A1(n24024), .A2(n25627), .B1(n24864), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_21/N3 ) );
  AOI22_X1 U13509 ( .A1(n24012), .A2(n25655), .B1(n25270), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_6/N3 ) );
  AOI22_X1 U13663 ( .A1(n24013), .A2(n25655), .B1(n25280), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_6/N3 ) );
  AOI22_X1 U13713 ( .A1(n24014), .A2(n26748), .B1(n25285), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_6/N3 ) );
  AOI22_X1 U13781 ( .A1(n23997), .A2(n25630), .B1(n25087), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_23/N3 ) );
  AOI22_X1 U13630 ( .A1(n24024), .A2(n25630), .B1(n24865), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_23/N3 ) );
  AOI22_X1 U13576 ( .A1(n24022), .A2(n26759), .B1(n24882), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_24/N3 ) );
  AOI22_X1 U13790 ( .A1(n23997), .A2(n25622), .B1(n25085), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_19/N3 ) );
  AOI22_X1 U13763 ( .A1(n23997), .A2(n25650), .B1(n2175), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_4/N3 ) );
  AOI22_X1 U13612 ( .A1(n24024), .A2(n25650), .B1(n2179), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_4/N3 ) );
  AOI22_X1 U13558 ( .A1(n24022), .A2(n26748), .B1(n2106), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_6/N3 ) );
  AOI22_X1 U13610 ( .A1(n24024), .A2(n25654), .B1(n2107), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_6/N3 ) );
  AOI22_X1 U13761 ( .A1(n23997), .A2(n25654), .B1(n2103), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_6/N3 ) );
  AOI22_X1 U13560 ( .A1(n24022), .A2(n26750), .B1(n2178), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_4/N3 ) );
  AOI22_X1 U13639 ( .A1(n24024), .A2(n25622), .B1(n24863), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_19/N3 ) );
  AOI22_X1 U13587 ( .A1(n24022), .A2(n26765), .B1(n24879), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_19/N3 ) );
  AOI22_X1 U13628 ( .A1(n24024), .A2(n25632), .B1(n24866), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_24/N3 ) );
  AOI22_X1 U13779 ( .A1(n23997), .A2(n25632), .B1(n25088), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_24/N3 ) );
  AOI22_X1 U13603 ( .A1(n24022), .A2(n26775), .B1(n3134), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_0/N3 ) );
  AOI22_X1 U13655 ( .A1(n24024), .A2(n25602), .B1(n3135), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_0/N3 ) );
  AOI22_X1 U13806 ( .A1(n23997), .A2(n25602), .B1(n3130), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_0/N3 ) );
  AOI22_X1 U13717 ( .A1(n24014), .A2(n26750), .B1(n24857), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_4/N3 ) );
  AOI22_X1 U13507 ( .A1(n24012), .A2(n25657), .B1(n24890), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_7/N3 ) );
  AOI22_X1 U13661 ( .A1(n24013), .A2(n25657), .B1(n24845), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_7/N3 ) );
  AOI22_X1 U13711 ( .A1(n24014), .A2(n26747), .B1(n25037), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_7/N3 ) );
  AOI22_X1 U13667 ( .A1(n24013), .A2(n25651), .B1(n25281), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_4/N3 ) );
  AOI22_X1 U13513 ( .A1(n24012), .A2(n25651), .B1(n25039), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_4/N3 ) );
  AOI22_X1 U13679 ( .A1(n24013), .A2(n25631), .B1(n774), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_23/N3 ) );
  AOI22_X1 U13735 ( .A1(n24014), .A2(n26765), .B1(n891), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_19/N3 ) );
  AOI22_X1 U13578 ( .A1(n24022), .A2(n26760), .B1(n24881), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_23/N3 ) );
  AOI22_X1 U13557 ( .A1(n24022), .A2(n26747), .B1(n2070), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_7/N3 ) );
  AOI22_X1 U13609 ( .A1(n24024), .A2(n25656), .B1(n2071), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_7/N3 ) );
  AOI22_X1 U13760 ( .A1(n23997), .A2(n25656), .B1(n2067), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_7/N3 ) );
  AOI22_X1 U13794 ( .A1(n23997), .A2(n25618), .B1(n25083), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_17/N3 ) );
  AOI22_X1 U13685 ( .A1(n24013), .A2(n25623), .B1(n892), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_19/N3 ) );
  AOI22_X1 U13532 ( .A1(n24012), .A2(n25623), .B1(n893), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_19/N3 ) );
  AOI22_X1 U13785 ( .A1(n23997), .A2(n25627), .B1(n25086), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_21/N3 ) );
  AOI22_X1 U13505 ( .A1(n24012), .A2(n25659), .B1(n24891), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_8/N3 ) );
  AOI22_X1 U13659 ( .A1(n24013), .A2(n25659), .B1(n24846), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_8/N3 ) );
  AOI22_X1 U13709 ( .A1(n24014), .A2(n26746), .B1(n25038), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_8/N3 ) );
  AOI22_X1 U13768 ( .A1(n23997), .A2(n25644), .B1(n2211), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_3/N3 ) );
  AOI22_X1 U13759 ( .A1(n23997), .A2(n25658), .B1(n2031), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_8/N3 ) );
  AOI22_X1 U13617 ( .A1(n24024), .A2(n25644), .B1(n2215), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_3/N3 ) );
  AOI22_X1 U13565 ( .A1(n24022), .A2(n26753), .B1(n2214), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_3/N3 ) );
  AOI22_X1 U13523 ( .A1(n24012), .A2(n25637), .B1(n620), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_26/N3 ) );
  AOI22_X1 U13548 ( .A1(n24012), .A2(n25605), .B1(n25099), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_1/N3 ) );
  AOI22_X1 U13792 ( .A1(n23997), .A2(n25620), .B1(n25084), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_18/N3 ) );
  AOI22_X1 U13641 ( .A1(n24024), .A2(n25620), .B1(n24862), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_18/N3 ) );
  AOI22_X1 U13701 ( .A1(n24013), .A2(n25605), .B1(n25272), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_1/N3 ) );
  AOI22_X1 U13751 ( .A1(n24014), .A2(n26774), .B1(n24851), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_1/N3 ) );
  AOI22_X1 U13527 ( .A1(n24012), .A2(n25629), .B1(n814), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_22/N3 ) );
  AOI22_X1 U13556 ( .A1(n24022), .A2(n26746), .B1(n2034), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_8/N3 ) );
  AOI22_X1 U13608 ( .A1(n24024), .A2(n25658), .B1(n2035), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_8/N3 ) );
  AOI22_X1 U13589 ( .A1(n24022), .A2(n26766), .B1(n24878), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_18/N3 ) );
  AOI22_X1 U13680 ( .A1(n24013), .A2(n25629), .B1(n813), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_22/N3 ) );
  AOI22_X1 U13533 ( .A1(n24012), .A2(n25621), .B1(n932), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_18/N3 ) );
  AOI22_X1 U13624 ( .A1(n24024), .A2(n25636), .B1(n24868), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_26/N3 ) );
  AOI22_X1 U13775 ( .A1(n23997), .A2(n25636), .B1(n25090), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_26/N3 ) );
  AOI22_X1 U13730 ( .A1(n24014), .A2(n26761), .B1(n812), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_22/N3 ) );
  AOI22_X1 U13676 ( .A1(n24013), .A2(n25637), .B1(n619), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_26/N3 ) );
  AOI22_X1 U13686 ( .A1(n24013), .A2(n25621), .B1(n931), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_18/N3 ) );
  AOI22_X1 U13726 ( .A1(n24014), .A2(n26757), .B1(n618), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_26/N3 ) );
  AOI22_X1 U13736 ( .A1(n24014), .A2(n26766), .B1(n930), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_18/N3 ) );
  AOI22_X1 U13729 ( .A1(n24014), .A2(n26760), .B1(n773), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_23/N3 ) );
  AOI22_X1 U13687 ( .A1(n24013), .A2(n25619), .B1(n698), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_17/N3 ) );
  AOI22_X1 U13572 ( .A1(n24022), .A2(n26757), .B1(n24884), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_26/N3 ) );
  AOI22_X1 U13563 ( .A1(n20611), .A2(n26752), .B1(n24888), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_30/N3 ) );
  AOI22_X1 U13725 ( .A1(n20667), .A2(n26756), .B1(n579), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_27/N3 ) );
  AOI22_X1 U13570 ( .A1(n20611), .A2(n26756), .B1(n24885), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_27/N3 ) );
  AOI22_X1 U13522 ( .A1(n20592), .A2(n25639), .B1(n581), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_27/N3 ) );
  AOI22_X1 U13670 ( .A1(n20650), .A2(n25647), .B1(n501), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_30/N3 ) );
  AOI22_X1 U13517 ( .A1(n20592), .A2(n25647), .B1(n502), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_30/N3 ) );
  AOI22_X1 U13766 ( .A1(n23997), .A2(n25646), .B1(n25094), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_30/N3 ) );
  AOI22_X1 U13675 ( .A1(n20650), .A2(n25639), .B1(n580), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_27/N3 ) );
  AOI22_X1 U13799 ( .A1(n23997), .A2(n25612), .B1(n2931), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_14/N3 ) );
  AOI22_X1 U13615 ( .A1(n20630), .A2(n25646), .B1(n24872), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_30/N3 ) );
  AOI22_X1 U13529 ( .A1(n20592), .A2(n25626), .B1(n854), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_20/N3 ) );
  AOI22_X1 U13773 ( .A1(n23997), .A2(n25638), .B1(n25091), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_27/N3 ) );
  AOI22_X1 U13682 ( .A1(n20650), .A2(n25626), .B1(n853), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_20/N3 ) );
  AOI22_X1 U13648 ( .A1(n20630), .A2(n25612), .B1(n2935), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_14/N3 ) );
  AOI22_X1 U13596 ( .A1(n20611), .A2(n26770), .B1(n2934), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_14/N3 ) );
  AOI22_X1 U13732 ( .A1(n20667), .A2(n26763), .B1(n852), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_20/N3 ) );
  AOI22_X1 U13787 ( .A1(n23997), .A2(net717157), .B1(net740972), .B2(n20686), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_10/DFF_20/N3 ) );
  AOI22_X1 U13636 ( .A1(n20630), .A2(net717157), .B1(net741216), .B2(n20632), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_13/DFF_20/N3 ) );
  AOI22_X1 U13584 ( .A1(n20611), .A2(n26763), .B1(net741198), .B2(n20613), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_14/DFF_20/N3 ) );
  AOI22_X1 U13720 ( .A1(n20667), .A2(n26752), .B1(n500), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_30/N3 ) );
  AOI22_X1 U13741 ( .A1(n20667), .A2(n26770), .B1(n24855), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_14/N3 ) );
  AOI22_X1 U13691 ( .A1(n20650), .A2(n25613), .B1(n25275), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_14/N3 ) );
  AOI22_X1 U13622 ( .A1(n20630), .A2(n25638), .B1(n24869), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_27/N3 ) );
  AOI22_X1 U13538 ( .A1(n20592), .A2(n25613), .B1(n25103), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_14/N3 ) );
  AOI22_X1 U13566 ( .A1(n20611), .A2(n26754), .B1(n24887), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_29/N3 ) );
  AOI22_X1 U13618 ( .A1(n20630), .A2(n25642), .B1(n24871), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_29/N3 ) );
  AOI22_X1 U13554 ( .A1(n20611), .A2(n26745), .B1(n25303), .B2(n20613), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_9/N3 ) );
  AOI22_X1 U13504 ( .A1(n20592), .A2(n25661), .B1(n352), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_9/N3 ) );
  AOI22_X1 U13673 ( .A1(n20650), .A2(n25643), .B1(n427), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_29/N3 ) );
  AOI22_X1 U13769 ( .A1(n23997), .A2(n25642), .B1(n25093), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_29/N3 ) );
  AOI22_X1 U13520 ( .A1(n20592), .A2(n25643), .B1(n428), .B2(n20593), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_29/N3 ) );
  AOI22_X1 U13606 ( .A1(n20630), .A2(n25660), .B1(n24874), .B2(n20632), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_9/N3 ) );
  AOI22_X1 U13757 ( .A1(n23997), .A2(n25660), .B1(n25096), .B2(n20686), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_9/N3 ) );
  AOI22_X1 U13658 ( .A1(n20650), .A2(n25661), .B1(n351), .B2(n20651), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_9/N3 ) );
  AOI22_X1 U13723 ( .A1(n20667), .A2(n26754), .B1(n426), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_29/N3 ) );
  AOI22_X1 U13708 ( .A1(n20667), .A2(n26745), .B1(n350), .B2(n20668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_9/N3 ) );
  AOI22_X1 U12978 ( .A1(n24002), .A2(net717153), .B1(net741518), .B2(n20394), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_24/DFF_22/N3 ) );
  AOI22_X1 U12927 ( .A1(n24003), .A2(n26761), .B1(net741108), .B2(n20375), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_25/DFF_22/N3 ) );
  AOI22_X1 U12991 ( .A1(n24002), .A2(n25616), .B1(n24641), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_16/N3 ) );
  AOI22_X1 U12963 ( .A1(n24002), .A2(n25644), .B1(n2196), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_3/N3 ) );
  AOI22_X1 U12998 ( .A1(n24002), .A2(n25606), .B1(n3060), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_10/N3 ) );
  AOI22_X1 U12548 ( .A1(n24025), .A2(n25651), .B1(n24777), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_4/N3 ) );
  AOI22_X1 U12629 ( .A1(n24018), .A2(n26761), .B1(net740858), .B2(n20296), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_30/DFF_22/N3 ) );
  AOI22_X1 U12947 ( .A1(n24003), .A2(n26773), .B1(n3059), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_10/N3 ) );
  AOI22_X1 U12865 ( .A1(n24009), .A2(n25645), .B1(n24650), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_3/N3 ) );
  AOI22_X1 U12649 ( .A1(n24018), .A2(n26773), .B1(n3062), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_10/N3 ) );
  AOI22_X1 U12579 ( .A1(n24025), .A2(n25621), .B1(n25210), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_18/N3 ) );
  AOI22_X1 U12912 ( .A1(n24003), .A2(n26753), .B1(n2195), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_3/N3 ) );
  AOI22_X1 U12763 ( .A1(n24004), .A2(n26750), .B1(n25080), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_4/N3 ) );
  AOI22_X1 U12642 ( .A1(n24018), .A2(n26768), .B1(n25186), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_16/N3 ) );
  AOI22_X1 U12989 ( .A1(n24002), .A2(n25618), .B1(n24642), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_17/N3 ) );
  AOI22_X1 U12714 ( .A1(n24006), .A2(n25651), .B1(n25044), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_4/N3 ) );
  AOI22_X1 U12893 ( .A1(n24009), .A2(n25607), .B1(n24632), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_10/N3 ) );
  AOI22_X1 U12844 ( .A1(n24005), .A2(n25606), .B1(n24631), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_10/N3 ) );
  AOI22_X1 U12795 ( .A1(n24004), .A2(n26773), .B1(n25177), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_10/N3 ) );
  AOI22_X1 U12609 ( .A1(n24018), .A2(n26750), .B1(n2162), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_4/N3 ) );
  AOI22_X1 U12874 ( .A1(n24009), .A2(n25629), .B1(n820), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_22/N3 ) );
  AOI22_X1 U12825 ( .A1(n24005), .A2(net717153), .B1(n821), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_22/N3 ) );
  AOI22_X1 U12638 ( .A1(n24018), .A2(n26766), .B1(n25188), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_18/N3 ) );
  AOI22_X1 U12970 ( .A1(n24002), .A2(n25636), .B1(n24625), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_26/N3 ) );
  AOI22_X1 U12614 ( .A1(n24018), .A2(n26753), .B1(n2198), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_3/N3 ) );
  AOI22_X1 U12936 ( .A1(n24003), .A2(n26766), .B1(n24958), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_18/N3 ) );
  AOI22_X1 U12987 ( .A1(n24002), .A2(n25620), .B1(n24622), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_18/N3 ) );
  AOI22_X1 U12919 ( .A1(n24003), .A2(n26757), .B1(n24964), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_26/N3 ) );
  AOI22_X1 U12621 ( .A1(n24018), .A2(n26757), .B1(n25194), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_26/N3 ) );
  AOI22_X1 U12746 ( .A1(n24006), .A2(n25607), .B1(n24973), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_10/N3 ) );
  AOI22_X1 U12595 ( .A1(n24025), .A2(n25607), .B1(n25203), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_10/N3 ) );
  AOI22_X1 U12733 ( .A1(n24006), .A2(n25621), .B1(n941), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_18/N3 ) );
  AOI22_X1 U12782 ( .A1(n24004), .A2(n26766), .B1(n940), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_18/N3 ) );
  AOI22_X1 U12831 ( .A1(n24005), .A2(n25620), .B1(n939), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_18/N3 ) );
  AOI22_X1 U12880 ( .A1(n24009), .A2(n25621), .B1(n938), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_18/N3 ) );
  AOI22_X1 U12954 ( .A1(n24002), .A2(n25658), .B1(n2016), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_8/N3 ) );
  AOI22_X1 U12903 ( .A1(n24003), .A2(n26746), .B1(n2015), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_8/N3 ) );
  AOI22_X1 U12605 ( .A1(n24018), .A2(n26746), .B1(n2018), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_8/N3 ) );
  AOI22_X1 U12812 ( .A1(n24005), .A2(n25650), .B1(n24775), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_4/N3 ) );
  AOI22_X1 U12861 ( .A1(n24009), .A2(n25651), .B1(n24776), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_4/N3 ) );
  AOI22_X1 U12940 ( .A1(n24003), .A2(n26768), .B1(n24956), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_16/N3 ) );
  AOI22_X1 U12853 ( .A1(n24009), .A2(n25659), .B1(n24664), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_8/N3 ) );
  AOI22_X1 U12804 ( .A1(n24005), .A2(n25658), .B1(n24665), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_8/N3 ) );
  AOI22_X1 U12776 ( .A1(n24004), .A2(n26761), .B1(n822), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_22/N3 ) );
  AOI22_X1 U12823 ( .A1(n24005), .A2(n25632), .B1(n667), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_24/N3 ) );
  AOI22_X1 U12727 ( .A1(n24006), .A2(n25629), .B1(n823), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_22/N3 ) );
  AOI22_X1 U12577 ( .A1(n24025), .A2(n25623), .B1(n25211), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_19/N3 ) );
  AOI22_X1 U12732 ( .A1(n24006), .A2(n25623), .B1(n902), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_19/N3 ) );
  AOI22_X1 U12781 ( .A1(n24004), .A2(n26765), .B1(n901), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_19/N3 ) );
  AOI22_X1 U12830 ( .A1(n24005), .A2(n25622), .B1(n900), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_19/N3 ) );
  AOI22_X1 U12879 ( .A1(n24009), .A2(n25623), .B1(n899), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_19/N3 ) );
  AOI22_X1 U12569 ( .A1(n24025), .A2(n25629), .B1(net740834), .B2(n20263), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_31/DFF_22/N3 ) );
  AOI22_X1 U12565 ( .A1(n24025), .A2(n25633), .B1(n25214), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_24/N3 ) );
  AOI22_X1 U12725 ( .A1(n24006), .A2(n25633), .B1(n669), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_24/N3 ) );
  AOI22_X1 U12870 ( .A1(n24009), .A2(n25637), .B1(n626), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_26/N3 ) );
  AOI22_X1 U12821 ( .A1(n24005), .A2(n25636), .B1(n627), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_26/N3 ) );
  AOI22_X1 U12755 ( .A1(n24004), .A2(n26746), .B1(n25185), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_8/N3 ) );
  AOI22_X1 U12706 ( .A1(n24006), .A2(n25659), .B1(n24983), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_8/N3 ) );
  AOI22_X1 U12540 ( .A1(n24025), .A2(n25659), .B1(n25049), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_8/N3 ) );
  AOI22_X1 U12772 ( .A1(n24004), .A2(n26757), .B1(n628), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_26/N3 ) );
  AOI22_X1 U12723 ( .A1(n24006), .A2(n25637), .B1(n629), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_26/N3 ) );
  AOI22_X1 U12561 ( .A1(n24025), .A2(n25637), .B1(n25216), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_26/N3 ) );
  AOI22_X1 U12955 ( .A1(n24002), .A2(n25656), .B1(n2052), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_7/N3 ) );
  AOI22_X1 U12636 ( .A1(n24018), .A2(n26765), .B1(n25189), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_19/N3 ) );
  AOI22_X1 U12904 ( .A1(n24003), .A2(n26747), .B1(n2051), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_7/N3 ) );
  AOI22_X1 U12934 ( .A1(n24003), .A2(n26765), .B1(n24959), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_19/N3 ) );
  AOI22_X1 U12985 ( .A1(n24002), .A2(n25622), .B1(n24643), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_19/N3 ) );
  AOI22_X1 U12606 ( .A1(n24018), .A2(n26747), .B1(n2054), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_7/N3 ) );
  AOI22_X1 U12550 ( .A1(n24025), .A2(n25649), .B1(n1755), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_31/N3 ) );
  AOI22_X1 U12855 ( .A1(n24009), .A2(n25657), .B1(n24660), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_7/N3 ) );
  AOI22_X1 U12806 ( .A1(n24005), .A2(n25656), .B1(n24661), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_7/N3 ) );
  AOI22_X1 U12757 ( .A1(n24004), .A2(n26747), .B1(n25184), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_7/N3 ) );
  AOI22_X1 U12708 ( .A1(n24006), .A2(n25657), .B1(n24982), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_7/N3 ) );
  AOI22_X1 U12542 ( .A1(n24025), .A2(n25657), .B1(n25048), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_7/N3 ) );
  AOI22_X1 U12956 ( .A1(n24002), .A2(n25654), .B1(n2088), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_6/N3 ) );
  AOI22_X1 U12905 ( .A1(n24003), .A2(n26748), .B1(n2087), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_6/N3 ) );
  AOI22_X1 U12607 ( .A1(n24018), .A2(n26748), .B1(n2090), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_6/N3 ) );
  AOI22_X1 U12857 ( .A1(n24009), .A2(n25655), .B1(n24672), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_6/N3 ) );
  AOI22_X1 U12808 ( .A1(n24005), .A2(n25654), .B1(n24658), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_6/N3 ) );
  AOI22_X1 U12907 ( .A1(n24003), .A2(n26750), .B1(n2159), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_4/N3 ) );
  AOI22_X1 U12958 ( .A1(n24002), .A2(n25650), .B1(n2160), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_4/N3 ) );
  AOI22_X1 U12546 ( .A1(n24025), .A2(n25653), .B1(n25277), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_5/N3 ) );
  AOI22_X1 U12712 ( .A1(n24006), .A2(n25653), .B1(n24980), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_5/N3 ) );
  AOI22_X1 U12774 ( .A1(n24004), .A2(n26759), .B1(n668), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_24/N3 ) );
  AOI22_X1 U12761 ( .A1(n24004), .A2(n26749), .B1(n25183), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_5/N3 ) );
  AOI22_X1 U12810 ( .A1(n24005), .A2(n25652), .B1(n24657), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_5/N3 ) );
  AOI22_X1 U12859 ( .A1(n24009), .A2(n25653), .B1(n24669), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_5/N3 ) );
  AOI22_X1 U12974 ( .A1(n24002), .A2(n25632), .B1(n24645), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_24/N3 ) );
  AOI22_X1 U12923 ( .A1(n24003), .A2(n26759), .B1(n24962), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_24/N3 ) );
  AOI22_X1 U12625 ( .A1(n24018), .A2(n26759), .B1(n25192), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_24/N3 ) );
  AOI22_X1 U12759 ( .A1(n24004), .A2(n26748), .B1(n25287), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_6/N3 ) );
  AOI22_X1 U12710 ( .A1(n24006), .A2(n25655), .B1(n24981), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_6/N3 ) );
  AOI22_X1 U12544 ( .A1(n24025), .A2(n25655), .B1(n25278), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_6/N3 ) );
  AOI22_X1 U12957 ( .A1(n24002), .A2(n25652), .B1(n2124), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_5/N3 ) );
  AOI22_X1 U12906 ( .A1(n24003), .A2(n26749), .B1(n2123), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_5/N3 ) );
  AOI22_X1 U12608 ( .A1(n24018), .A2(n26749), .B1(n2126), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_5/N3 ) );
  AOI22_X1 U12785 ( .A1(n24004), .A2(n26769), .B1(n25181), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_15/N3 ) );
  AOI22_X1 U12750 ( .A1(n24006), .A2(n25603), .B1(n24971), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_0/N3 ) );
  AOI22_X1 U12799 ( .A1(n24004), .A2(n26775), .B1(n25175), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_0/N3 ) );
  AOI22_X1 U12863 ( .A1(n24009), .A2(n25649), .B1(n470), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_31/N3 ) );
  AOI22_X1 U12814 ( .A1(n24005), .A2(n25648), .B1(n471), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_31/N3 ) );
  AOI22_X1 U12765 ( .A1(n24004), .A2(n26751), .B1(n472), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_31/N3 ) );
  AOI22_X1 U12631 ( .A1(n24018), .A2(n26762), .B1(n25190), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_21/N3 ) );
  AOI22_X1 U12716 ( .A1(n24006), .A2(n25649), .B1(n473), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_31/N3 ) );
  AOI22_X1 U12929 ( .A1(n24003), .A2(n26762), .B1(n24960), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_21/N3 ) );
  AOI22_X1 U12980 ( .A1(n24002), .A2(n25627), .B1(n24624), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_21/N3 ) );
  AOI22_X1 U12875 ( .A1(n24009), .A2(n25628), .B1(n743), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_21/N3 ) );
  AOI22_X1 U12826 ( .A1(n24005), .A2(n25627), .B1(n744), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_21/N3 ) );
  AOI22_X1 U12777 ( .A1(n24004), .A2(n26762), .B1(n745), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_21/N3 ) );
  AOI22_X1 U12728 ( .A1(n24006), .A2(n25628), .B1(n746), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_21/N3 ) );
  AOI22_X1 U12571 ( .A1(n24025), .A2(n25628), .B1(n25212), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_21/N3 ) );
  AOI22_X1 U12848 ( .A1(n24005), .A2(n25602), .B1(n24627), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_0/N3 ) );
  AOI22_X1 U12897 ( .A1(n24009), .A2(n25603), .B1(n24628), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_0/N3 ) );
  AOI22_X1 U12610 ( .A1(n24018), .A2(n26751), .B1(n25199), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_31/N3 ) );
  AOI22_X1 U12908 ( .A1(n24003), .A2(n26751), .B1(n24969), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_31/N3 ) );
  AOI22_X1 U12959 ( .A1(n24002), .A2(n25648), .B1(n24954), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_31/N3 ) );
  AOI22_X1 U12651 ( .A1(n24018), .A2(n26775), .B1(n3107), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_0/N3 ) );
  AOI22_X1 U12949 ( .A1(n24003), .A2(n26775), .B1(n3102), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_0/N3 ) );
  AOI22_X1 U13000 ( .A1(n24002), .A2(n25602), .B1(n3103), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_0/N3 ) );
  AOI22_X1 U12597 ( .A1(n24025), .A2(n25605), .B1(n25202), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_1/N3 ) );
  AOI22_X1 U12585 ( .A1(n24025), .A2(n25615), .B1(n25207), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_15/N3 ) );
  AOI22_X1 U12736 ( .A1(n24006), .A2(n25615), .B1(n24977), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_15/N3 ) );
  AOI22_X1 U12599 ( .A1(n24025), .A2(n25603), .B1(n25201), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_0/N3 ) );
  AOI22_X1 U12834 ( .A1(n24005), .A2(n25614), .B1(n24639), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_15/N3 ) );
  AOI22_X1 U12883 ( .A1(n24009), .A2(n25615), .B1(n24640), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_15/N3 ) );
  AOI22_X1 U12748 ( .A1(n24006), .A2(n25605), .B1(n24972), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_1/N3 ) );
  AOI22_X1 U12797 ( .A1(n24004), .A2(n26774), .B1(n25176), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_1/N3 ) );
  AOI22_X1 U12846 ( .A1(n24005), .A2(n25604), .B1(n24629), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_1/N3 ) );
  AOI22_X1 U12895 ( .A1(n24009), .A2(n25605), .B1(n24630), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_1/N3 ) );
  AOI22_X1 U12650 ( .A1(n24018), .A2(n26774), .B1(n2702), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_1/N3 ) );
  AOI22_X1 U12976 ( .A1(n24002), .A2(n25630), .B1(n24644), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_23/N3 ) );
  AOI22_X1 U12925 ( .A1(n24003), .A2(n26760), .B1(n24961), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_23/N3 ) );
  AOI22_X1 U12948 ( .A1(n24003), .A2(n26774), .B1(n2699), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_1/N3 ) );
  AOI22_X1 U12627 ( .A1(n24018), .A2(n26760), .B1(n25191), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_23/N3 ) );
  AOI22_X1 U12581 ( .A1(n24025), .A2(n25619), .B1(n25209), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_17/N3 ) );
  AOI22_X1 U12734 ( .A1(n24006), .A2(n25619), .B1(n708), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_17/N3 ) );
  AOI22_X1 U12644 ( .A1(n24018), .A2(n26769), .B1(n2882), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_15/N3 ) );
  AOI22_X1 U12783 ( .A1(n24004), .A2(n26767), .B1(n707), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_17/N3 ) );
  AOI22_X1 U12942 ( .A1(n24003), .A2(n26769), .B1(n2879), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_15/N3 ) );
  AOI22_X1 U12993 ( .A1(n24002), .A2(n25614), .B1(n2880), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_15/N3 ) );
  AOI22_X1 U12832 ( .A1(n24005), .A2(n25618), .B1(n706), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_17/N3 ) );
  AOI22_X1 U12999 ( .A1(n24002), .A2(n25604), .B1(n2700), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_1/N3 ) );
  AOI22_X1 U12575 ( .A1(n24025), .A2(n25625), .B1(n25304), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_2/N3 ) );
  AOI22_X1 U12563 ( .A1(n24025), .A2(n25635), .B1(n25215), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_25/N3 ) );
  AOI22_X1 U12724 ( .A1(n24006), .A2(n25635), .B1(n399), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_25/N3 ) );
  AOI22_X1 U12773 ( .A1(n24004), .A2(n26758), .B1(n398), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_25/N3 ) );
  AOI22_X1 U12730 ( .A1(n24006), .A2(n25625), .B1(n24978), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_2/N3 ) );
  AOI22_X1 U12938 ( .A1(n24003), .A2(n26767), .B1(n24957), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_17/N3 ) );
  AOI22_X1 U12881 ( .A1(n24009), .A2(n25619), .B1(n705), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_17/N3 ) );
  AOI22_X1 U12589 ( .A1(n24025), .A2(n25611), .B1(n25205), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_13/N3 ) );
  AOI22_X1 U12740 ( .A1(n24006), .A2(n25611), .B1(n24975), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_13/N3 ) );
  AOI22_X1 U12789 ( .A1(n24004), .A2(n26771), .B1(n25179), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_13/N3 ) );
  AOI22_X1 U12838 ( .A1(n24005), .A2(n25610), .B1(n25174), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_13/N3 ) );
  AOI22_X1 U12887 ( .A1(n24009), .A2(n25611), .B1(n24635), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_13/N3 ) );
  AOI22_X1 U12873 ( .A1(n24009), .A2(n25631), .B1(n781), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_23/N3 ) );
  AOI22_X1 U12966 ( .A1(n24002), .A2(n25640), .B1(n24648), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_28/N3 ) );
  AOI22_X1 U12915 ( .A1(n24003), .A2(n26755), .B1(n24966), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_28/N3 ) );
  AOI22_X1 U12617 ( .A1(n24018), .A2(n26755), .B1(n25196), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_28/N3 ) );
  AOI22_X1 U12822 ( .A1(n24005), .A2(n25634), .B1(n397), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_25/N3 ) );
  AOI22_X1 U12871 ( .A1(n24009), .A2(n25635), .B1(n396), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_25/N3 ) );
  AOI22_X1 U12824 ( .A1(n24005), .A2(n25630), .B1(n782), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_23/N3 ) );
  AOI22_X1 U12775 ( .A1(n24004), .A2(n26760), .B1(n783), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_23/N3 ) );
  AOI22_X1 U12726 ( .A1(n24006), .A2(n25631), .B1(n784), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_23/N3 ) );
  AOI22_X1 U12567 ( .A1(n24025), .A2(n25631), .B1(n25213), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_23/N3 ) );
  AOI22_X1 U12779 ( .A1(n24004), .A2(n26764), .B1(n25286), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_2/N3 ) );
  AOI22_X1 U12828 ( .A1(n24005), .A2(n25624), .B1(n24623), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_2/N3 ) );
  AOI22_X1 U12646 ( .A1(n24018), .A2(n26771), .B1(n2954), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_13/N3 ) );
  AOI22_X1 U12877 ( .A1(n24009), .A2(n25625), .B1(n24675), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_2/N3 ) );
  AOI22_X1 U12944 ( .A1(n24003), .A2(n26771), .B1(n2951), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_13/N3 ) );
  AOI22_X1 U12995 ( .A1(n24002), .A2(n25610), .B1(n2952), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_13/N3 ) );
  AOI22_X1 U12635 ( .A1(n24018), .A2(n26764), .B1(n2306), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_2/N3 ) );
  AOI22_X1 U12933 ( .A1(n24003), .A2(n26764), .B1(n2303), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_2/N3 ) );
  AOI22_X1 U12868 ( .A1(n24009), .A2(n25641), .B1(n548), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_28/N3 ) );
  AOI22_X1 U12819 ( .A1(n24005), .A2(n25640), .B1(n549), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_28/N3 ) );
  AOI22_X1 U12997 ( .A1(n24002), .A2(n25608), .B1(n3024), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_11/N3 ) );
  AOI22_X1 U12946 ( .A1(n24003), .A2(n26772), .B1(n3023), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_11/N3 ) );
  AOI22_X1 U12984 ( .A1(n24002), .A2(n25624), .B1(n2304), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_2/N3 ) );
  AOI22_X1 U12770 ( .A1(n24004), .A2(n26755), .B1(n550), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_28/N3 ) );
  AOI22_X1 U12648 ( .A1(n24018), .A2(n26772), .B1(n3026), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_11/N3 ) );
  AOI22_X1 U12721 ( .A1(n24006), .A2(n25641), .B1(n551), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_28/N3 ) );
  AOI22_X1 U12623 ( .A1(n24018), .A2(n26758), .B1(n25193), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_25/N3 ) );
  AOI22_X1 U12557 ( .A1(n24025), .A2(n25641), .B1(n25218), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_28/N3 ) );
  AOI22_X1 U12921 ( .A1(n24003), .A2(n26758), .B1(n24963), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_25/N3 ) );
  AOI22_X1 U12583 ( .A1(n24025), .A2(n25617), .B1(n25208), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_16/N3 ) );
  AOI22_X1 U12735 ( .A1(n24006), .A2(n25617), .B1(n981), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_16/N3 ) );
  AOI22_X1 U12784 ( .A1(n24004), .A2(n26768), .B1(n980), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_16/N3 ) );
  AOI22_X1 U12833 ( .A1(n24005), .A2(n25616), .B1(n979), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_16/N3 ) );
  AOI22_X1 U12882 ( .A1(n24009), .A2(n25617), .B1(n978), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_16/N3 ) );
  AOI22_X1 U12972 ( .A1(n24002), .A2(n25634), .B1(n24646), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_25/N3 ) );
  AOI22_X1 U12553 ( .A1(n24025), .A2(n25645), .B1(n25047), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_3/N3 ) );
  AOI22_X1 U12718 ( .A1(n24006), .A2(n25645), .B1(n24979), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_3/N3 ) );
  AOI22_X1 U12767 ( .A1(n24004), .A2(n26753), .B1(n25182), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_3/N3 ) );
  AOI22_X1 U12891 ( .A1(n24009), .A2(n25609), .B1(n24634), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_11/N3 ) );
  AOI22_X1 U12842 ( .A1(n24005), .A2(n25608), .B1(n24633), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_11/N3 ) );
  AOI22_X1 U12793 ( .A1(n24004), .A2(n26772), .B1(n25178), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_11/N3 ) );
  AOI22_X1 U12744 ( .A1(n24006), .A2(n25609), .B1(n24974), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_11/N3 ) );
  AOI22_X1 U12593 ( .A1(n24025), .A2(n25609), .B1(n25204), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_11/N3 ) );
  AOI22_X1 U12816 ( .A1(n24005), .A2(n25644), .B1(n24651), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_3/N3 ) );
  AOI22_X1 U12640 ( .A1(n24018), .A2(n26767), .B1(n25187), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_17/N3 ) );
  AOI22_X1 U12872 ( .A1(n24009), .A2(n25633), .B1(n666), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_24/N3 ) );
  AOI22_X1 U12982 ( .A1(n24002), .A2(net717157), .B1(net741520), .B2(n20394), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_24/DFF_20/N3 ) );
  AOI22_X1 U12766 ( .A1(n24004), .A2(n26752), .B1(n510), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_30/N3 ) );
  AOI22_X1 U12931 ( .A1(n24003), .A2(n26763), .B1(net741110), .B2(n20375), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_25/DFF_20/N3 ) );
  AOI22_X1 U12885 ( .A1(n20370), .A2(n25613), .B1(n24638), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_14/N3 ) );
  AOI22_X1 U12913 ( .A1(n24003), .A2(n26754), .B1(n24967), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_29/N3 ) );
  AOI22_X1 U12615 ( .A1(n20294), .A2(n26754), .B1(n25197), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_29/N3 ) );
  AOI22_X1 U12633 ( .A1(n20294), .A2(n26763), .B1(net740860), .B2(n20296), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_30/DFF_20/N3 ) );
  AOI22_X1 U12901 ( .A1(n24003), .A2(n26745), .B1(n24970), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_9/N3 ) );
  AOI22_X1 U12994 ( .A1(n24002), .A2(n25612), .B1(n2916), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_14/N3 ) );
  AOI22_X1 U12943 ( .A1(n24003), .A2(n26770), .B1(n2915), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_14/N3 ) );
  AOI22_X1 U12876 ( .A1(n20370), .A2(n25626), .B1(n860), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_20/N3 ) );
  AOI22_X1 U12827 ( .A1(n24005), .A2(net717157), .B1(n861), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_20/N3 ) );
  AOI22_X1 U12778 ( .A1(n24004), .A2(n26763), .B1(n862), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_20/N3 ) );
  AOI22_X1 U12729 ( .A1(n24006), .A2(n25626), .B1(n863), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_20/N3 ) );
  AOI22_X1 U12573 ( .A1(n20261), .A2(n25626), .B1(net740836), .B2(n20263), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_31/DFF_20/N3 ) );
  AOI22_X1 U12555 ( .A1(n20261), .A2(n25643), .B1(n25219), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_29/N3 ) );
  AOI22_X1 U12754 ( .A1(n24004), .A2(n26745), .B1(n360), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_9/N3 ) );
  AOI22_X1 U12910 ( .A1(n24003), .A2(n26752), .B1(n24968), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_30/N3 ) );
  AOI22_X1 U12820 ( .A1(n24005), .A2(n25638), .B1(n588), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_27/N3 ) );
  AOI22_X1 U12869 ( .A1(n20370), .A2(n25639), .B1(n587), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_27/N3 ) );
  AOI22_X1 U12705 ( .A1(n24006), .A2(n25661), .B1(n361), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_9/N3 ) );
  AOI22_X1 U12538 ( .A1(n20261), .A2(n25661), .B1(n25221), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_9/N3 ) );
  AOI22_X1 U12964 ( .A1(n24002), .A2(n25642), .B1(n24626), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_29/N3 ) );
  AOI22_X1 U12917 ( .A1(n24003), .A2(n26756), .B1(n24965), .B2(n20375), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_27/N3 ) );
  AOI22_X1 U12968 ( .A1(n24002), .A2(n25638), .B1(n24647), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_27/N3 ) );
  AOI22_X1 U12952 ( .A1(n24002), .A2(n25660), .B1(n24955), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_9/N3 ) );
  AOI22_X1 U12836 ( .A1(n24005), .A2(n25612), .B1(n24637), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_14/N3 ) );
  AOI22_X1 U12603 ( .A1(n20294), .A2(n26745), .B1(n25200), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_9/N3 ) );
  AOI22_X1 U12559 ( .A1(n20261), .A2(n25639), .B1(n25217), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_27/N3 ) );
  AOI22_X1 U12722 ( .A1(n24006), .A2(n25639), .B1(n590), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_27/N3 ) );
  AOI22_X1 U12852 ( .A1(n20370), .A2(n25661), .B1(n358), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_9/N3 ) );
  AOI22_X1 U12803 ( .A1(n24005), .A2(n25660), .B1(n359), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_9/N3 ) );
  AOI22_X1 U12771 ( .A1(n24004), .A2(n26756), .B1(n589), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_27/N3 ) );
  AOI22_X1 U12720 ( .A1(n24006), .A2(n25643), .B1(n437), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_29/N3 ) );
  AOI22_X1 U12645 ( .A1(n20294), .A2(n26770), .B1(n2918), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_14/N3 ) );
  AOI22_X1 U12867 ( .A1(n20370), .A2(n25643), .B1(n434), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_29/N3 ) );
  AOI22_X1 U12818 ( .A1(n24005), .A2(n25642), .B1(n435), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_29/N3 ) );
  AOI22_X1 U12769 ( .A1(n24004), .A2(n26754), .B1(n436), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_29/N3 ) );
  AOI22_X1 U12587 ( .A1(n20261), .A2(n25613), .B1(n25206), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_14/N3 ) );
  AOI22_X1 U12961 ( .A1(n24002), .A2(n25646), .B1(n24653), .B2(n20394), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_30/N3 ) );
  AOI22_X1 U12612 ( .A1(n20294), .A2(n26752), .B1(n25198), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_30/N3 ) );
  AOI22_X1 U12619 ( .A1(n20294), .A2(n26756), .B1(n25195), .B2(n20296), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_27/N3 ) );
  AOI22_X1 U12864 ( .A1(n20370), .A2(n25647), .B1(n508), .B2(n20371), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_30/N3 ) );
  AOI22_X1 U12551 ( .A1(n20261), .A2(n25647), .B1(n25220), .B2(n20263), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_30/N3 ) );
  AOI22_X1 U12787 ( .A1(n24004), .A2(n26770), .B1(n25180), .B2(n20351), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_14/N3 ) );
  AOI22_X1 U12738 ( .A1(n24006), .A2(n25613), .B1(n24976), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_14/N3 ) );
  AOI22_X1 U12815 ( .A1(n24005), .A2(n25646), .B1(n509), .B2(n20368), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_30/N3 ) );
  AOI22_X1 U12717 ( .A1(n24006), .A2(n25647), .B1(n511), .B2(n20334), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_30/N3 ) );
  AOI22_X1 U13414 ( .A1(n23999), .A2(n26757), .B1(n24908), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_26/N3 ) );
  AOI22_X1 U13030 ( .A1(n24010), .A2(n25633), .B1(n25166), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_24/N3 ) );
  AOI22_X1 U13474 ( .A1(n23998), .A2(n25634), .B1(n391), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_25/N3 ) );
  AOI22_X1 U13475 ( .A1(n23998), .A2(n25632), .B1(n661), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_24/N3 ) );
  AOI22_X1 U13348 ( .A1(n24000), .A2(n25637), .B1(n25122), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_26/N3 ) );
  AOI22_X1 U13418 ( .A1(n23999), .A2(n26759), .B1(n24906), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_24/N3 ) );
  AOI22_X1 U13294 ( .A1(n23996), .A2(n25632), .B1(n25071), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_24/N3 ) );
  AOI22_X1 U13026 ( .A1(n24010), .A2(n25637), .B1(n25168), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_26/N3 ) );
  AOI22_X1 U13086 ( .A1(n24011), .A2(n26757), .B1(n624), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_26/N3 ) );
  AOI22_X1 U13028 ( .A1(n24010), .A2(n25635), .B1(n25167), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_25/N3 ) );
  AOI22_X1 U13434 ( .A1(n23999), .A2(n26767), .B1(n24900), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_17/N3 ) );
  AOI22_X1 U13473 ( .A1(n23998), .A2(n25636), .B1(n621), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_26/N3 ) );
  AOI22_X1 U13097 ( .A1(n24011), .A2(n26767), .B1(n703), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_17/N3 ) );
  AOI22_X1 U13088 ( .A1(n24011), .A2(n26759), .B1(n664), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_24/N3 ) );
  AOI22_X1 U13131 ( .A1(n24001), .A2(n25640), .B1(n24946), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_28/N3 ) );
  AOI22_X1 U13182 ( .A1(n24020), .A2(n25641), .B1(n25140), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_28/N3 ) );
  AOI22_X1 U13286 ( .A1(n23996), .A2(n25640), .B1(n25075), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_28/N3 ) );
  AOI22_X1 U13352 ( .A1(n24000), .A2(n25633), .B1(n25120), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_24/N3 ) );
  AOI22_X1 U13186 ( .A1(n24020), .A2(n25637), .B1(n25138), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_26/N3 ) );
  AOI22_X1 U13022 ( .A1(n24010), .A2(n25641), .B1(n25170), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_28/N3 ) );
  AOI22_X1 U13084 ( .A1(n24011), .A2(n26755), .B1(n546), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_28/N3 ) );
  AOI22_X1 U13344 ( .A1(n24000), .A2(n25641), .B1(n25124), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_28/N3 ) );
  AOI22_X1 U13079 ( .A1(n24011), .A2(n26751), .B1(n468), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_31/N3 ) );
  AOI22_X1 U13139 ( .A1(n24001), .A2(n25632), .B1(n24942), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_24/N3 ) );
  AOI22_X1 U13190 ( .A1(n24020), .A2(n25633), .B1(n25136), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_24/N3 ) );
  AOI22_X1 U13416 ( .A1(n23999), .A2(n26758), .B1(n24907), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_25/N3 ) );
  AOI22_X1 U13350 ( .A1(n24000), .A2(n25635), .B1(n25121), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_25/N3 ) );
  AOI22_X1 U13087 ( .A1(n24011), .A2(n26758), .B1(n394), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_25/N3 ) );
  AOI22_X1 U13309 ( .A1(n23996), .A2(n25618), .B1(n25066), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_17/N3 ) );
  AOI22_X1 U13205 ( .A1(n24020), .A2(n25619), .B1(n25131), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_17/N3 ) );
  AOI22_X1 U13368 ( .A1(n24000), .A2(n25619), .B1(n25115), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_17/N3 ) );
  AOI22_X1 U13154 ( .A1(n24001), .A2(n25618), .B1(n24937), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_17/N3 ) );
  AOI22_X1 U13046 ( .A1(n24010), .A2(n25619), .B1(n25161), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_17/N3 ) );
  AOI22_X1 U13279 ( .A1(n23996), .A2(n25648), .B1(n24654), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_31/N3 ) );
  AOI22_X1 U13175 ( .A1(n24020), .A2(n25649), .B1(n25143), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_31/N3 ) );
  AOI22_X1 U13124 ( .A1(n24001), .A2(n25648), .B1(n24949), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_31/N3 ) );
  AOI22_X1 U13135 ( .A1(n24001), .A2(n25636), .B1(n24944), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_26/N3 ) );
  AOI22_X1 U13300 ( .A1(n23996), .A2(n25627), .B1(n25069), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_21/N3 ) );
  AOI22_X1 U13290 ( .A1(n23996), .A2(n25636), .B1(n25073), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_26/N3 ) );
  AOI22_X1 U13292 ( .A1(n23996), .A2(n25634), .B1(n25072), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_25/N3 ) );
  AOI22_X1 U13188 ( .A1(n24020), .A2(n25635), .B1(n25137), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_25/N3 ) );
  AOI22_X1 U13137 ( .A1(n24001), .A2(n25634), .B1(n24943), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_25/N3 ) );
  AOI22_X1 U13467 ( .A1(n23998), .A2(n25648), .B1(n465), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_31/N3 ) );
  AOI22_X1 U13196 ( .A1(n24020), .A2(n25628), .B1(n25134), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_21/N3 ) );
  AOI22_X1 U13145 ( .A1(n24001), .A2(n25627), .B1(n24940), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_21/N3 ) );
  AOI22_X1 U13402 ( .A1(n23999), .A2(n26751), .B1(n24914), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_31/N3 ) );
  AOI22_X1 U13410 ( .A1(n23999), .A2(n26755), .B1(n24910), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_28/N3 ) );
  AOI22_X1 U13483 ( .A1(n23998), .A2(n25618), .B1(n700), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_17/N3 ) );
  AOI22_X1 U13471 ( .A1(n23998), .A2(n25640), .B1(n543), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_28/N3 ) );
  AOI22_X1 U13015 ( .A1(n24010), .A2(n25649), .B1(n469), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_31/N3 ) );
  AOI22_X1 U13336 ( .A1(n24000), .A2(n25649), .B1(n25127), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_31/N3 ) );
  AOI22_X1 U13328 ( .A1(n24000), .A2(n25657), .B1(n24589), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_7/N3 ) );
  AOI22_X1 U13485 ( .A1(n23998), .A2(n25614), .B1(n25268), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_15/N3 ) );
  AOI22_X1 U13372 ( .A1(n24000), .A2(n25615), .B1(n25113), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_15/N3 ) );
  AOI22_X1 U13077 ( .A1(n24011), .A2(n26750), .B1(n25152), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_4/N3 ) );
  AOI22_X1 U13099 ( .A1(n24011), .A2(n26769), .B1(n25151), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_15/N3 ) );
  AOI22_X1 U13050 ( .A1(n24010), .A2(n25615), .B1(n25159), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_15/N3 ) );
  AOI22_X1 U13013 ( .A1(n24010), .A2(n25651), .B1(n25041), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_4/N3 ) );
  AOI22_X1 U13158 ( .A1(n24001), .A2(n25614), .B1(n2876), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_15/N3 ) );
  AOI22_X1 U13209 ( .A1(n24020), .A2(n25615), .B1(n2877), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_15/N3 ) );
  AOI22_X1 U13283 ( .A1(n23996), .A2(n25644), .B1(n2190), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_3/N3 ) );
  AOI22_X1 U13313 ( .A1(n23996), .A2(n25614), .B1(n2874), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_15/N3 ) );
  AOI22_X1 U13179 ( .A1(n24020), .A2(n25645), .B1(n2193), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_3/N3 ) );
  AOI22_X1 U13128 ( .A1(n24001), .A2(n25644), .B1(n2192), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_3/N3 ) );
  AOI22_X1 U13334 ( .A1(n24000), .A2(n25651), .B1(n25128), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_4/N3 ) );
  AOI22_X1 U13400 ( .A1(n23999), .A2(n26750), .B1(n24915), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_4/N3 ) );
  AOI22_X1 U13465 ( .A1(n23998), .A2(n25650), .B1(n25326), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_4/N3 ) );
  AOI22_X1 U13054 ( .A1(n24010), .A2(n25611), .B1(n25157), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_13/N3 ) );
  AOI22_X1 U13103 ( .A1(n24011), .A2(n26771), .B1(n25149), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_13/N3 ) );
  AOI22_X1 U13376 ( .A1(n24000), .A2(n25611), .B1(n25111), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_13/N3 ) );
  AOI22_X1 U13442 ( .A1(n23999), .A2(n26771), .B1(n24896), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_13/N3 ) );
  AOI22_X1 U13489 ( .A1(n23998), .A2(n25610), .B1(n25305), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_13/N3 ) );
  AOI22_X1 U13160 ( .A1(n24001), .A2(n25610), .B1(n2948), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_13/N3 ) );
  AOI22_X1 U13211 ( .A1(n24020), .A2(n25611), .B1(n24636), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_13/N3 ) );
  AOI22_X1 U13469 ( .A1(n23998), .A2(n25644), .B1(n1442), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_3/N3 ) );
  AOI22_X1 U13315 ( .A1(n23996), .A2(n25610), .B1(n25046), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_13/N3 ) );
  AOI22_X1 U13406 ( .A1(n23999), .A2(n26753), .B1(n24912), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_3/N3 ) );
  AOI22_X1 U13340 ( .A1(n24000), .A2(n25645), .B1(n24588), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_3/N3 ) );
  AOI22_X1 U13123 ( .A1(n24001), .A2(n25650), .B1(n2156), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_4/N3 ) );
  AOI22_X1 U13081 ( .A1(n24011), .A2(n26753), .B1(n24652), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_3/N3 ) );
  AOI22_X1 U13018 ( .A1(n24010), .A2(n25645), .B1(n25040), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_3/N3 ) );
  AOI22_X1 U13048 ( .A1(n24010), .A2(n25617), .B1(n25160), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_16/N3 ) );
  AOI22_X1 U13098 ( .A1(n24011), .A2(n26768), .B1(n976), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_16/N3 ) );
  AOI22_X1 U13370 ( .A1(n24000), .A2(n25617), .B1(n25114), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_16/N3 ) );
  AOI22_X1 U13436 ( .A1(n23999), .A2(n26768), .B1(n24899), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_16/N3 ) );
  AOI22_X1 U13174 ( .A1(n24020), .A2(n25651), .B1(n2157), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_4/N3 ) );
  AOI22_X1 U13484 ( .A1(n23998), .A2(n25616), .B1(n973), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_16/N3 ) );
  AOI22_X1 U13278 ( .A1(n23996), .A2(n25650), .B1(n2154), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_4/N3 ) );
  AOI22_X1 U13011 ( .A1(n24010), .A2(n25653), .B1(n24952), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_5/N3 ) );
  AOI22_X1 U13304 ( .A1(n23996), .A2(n25624), .B1(n2298), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_2/N3 ) );
  AOI22_X1 U13075 ( .A1(n24011), .A2(n26749), .B1(n24670), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_5/N3 ) );
  AOI22_X1 U13200 ( .A1(n24020), .A2(n25625), .B1(n2301), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_2/N3 ) );
  AOI22_X1 U13149 ( .A1(n24001), .A2(n25624), .B1(n2300), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_2/N3 ) );
  AOI22_X1 U13156 ( .A1(n24001), .A2(n25616), .B1(n24936), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_16/N3 ) );
  AOI22_X1 U13207 ( .A1(n24020), .A2(n25617), .B1(n25130), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_16/N3 ) );
  AOI22_X1 U13311 ( .A1(n23996), .A2(n25616), .B1(n25065), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_16/N3 ) );
  AOI22_X1 U13332 ( .A1(n24000), .A2(n25653), .B1(n24592), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_5/N3 ) );
  AOI22_X1 U13044 ( .A1(n24010), .A2(n25621), .B1(n25162), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_18/N3 ) );
  AOI22_X1 U13398 ( .A1(n23999), .A2(n26749), .B1(n24916), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_5/N3 ) );
  AOI22_X1 U13096 ( .A1(n24011), .A2(n26766), .B1(n936), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_18/N3 ) );
  AOI22_X1 U13366 ( .A1(n24000), .A2(n25621), .B1(n25116), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_18/N3 ) );
  AOI22_X1 U13432 ( .A1(n23999), .A2(n26766), .B1(n24901), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_18/N3 ) );
  AOI22_X1 U13463 ( .A1(n23998), .A2(n25652), .B1(n25105), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_5/N3 ) );
  AOI22_X1 U13482 ( .A1(n23998), .A2(n25620), .B1(n933), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_18/N3 ) );
  AOI22_X1 U13318 ( .A1(n23996), .A2(n25608), .B1(n3018), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_11/N3 ) );
  AOI22_X1 U13214 ( .A1(n24020), .A2(n25609), .B1(n3021), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_11/N3 ) );
  AOI22_X1 U13480 ( .A1(n23998), .A2(n25624), .B1(n1481), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_2/N3 ) );
  AOI22_X1 U13162 ( .A1(n24001), .A2(n25608), .B1(n3020), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_11/N3 ) );
  AOI22_X1 U13428 ( .A1(n23999), .A2(n26764), .B1(n24903), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_2/N3 ) );
  AOI22_X1 U13152 ( .A1(n24001), .A2(n25620), .B1(n24938), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_18/N3 ) );
  AOI22_X1 U13203 ( .A1(n24020), .A2(n25621), .B1(n25132), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_18/N3 ) );
  AOI22_X1 U13362 ( .A1(n24000), .A2(n25625), .B1(n24676), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_2/N3 ) );
  AOI22_X1 U13093 ( .A1(n24011), .A2(n26764), .B1(n24594), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_2/N3 ) );
  AOI22_X1 U13122 ( .A1(n24001), .A2(n25652), .B1(n2120), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_5/N3 ) );
  AOI22_X1 U13493 ( .A1(n23998), .A2(n25608), .B1(n25266), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_11/N3 ) );
  AOI22_X1 U13307 ( .A1(n23996), .A2(n25620), .B1(n25067), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_18/N3 ) );
  AOI22_X1 U13040 ( .A1(n24010), .A2(n25625), .B1(n24951), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_2/N3 ) );
  AOI22_X1 U13446 ( .A1(n23999), .A2(n26772), .B1(n24895), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_11/N3 ) );
  AOI22_X1 U13380 ( .A1(n24000), .A2(n25609), .B1(n25110), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_11/N3 ) );
  AOI22_X1 U13042 ( .A1(n24010), .A2(n25623), .B1(n25163), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_19/N3 ) );
  AOI22_X1 U13095 ( .A1(n24011), .A2(n26765), .B1(n897), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_19/N3 ) );
  AOI22_X1 U13364 ( .A1(n24000), .A2(n25623), .B1(n25117), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_19/N3 ) );
  AOI22_X1 U13430 ( .A1(n23999), .A2(n26765), .B1(n24902), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_19/N3 ) );
  AOI22_X1 U13481 ( .A1(n23998), .A2(n25622), .B1(n894), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_19/N3 ) );
  AOI22_X1 U13173 ( .A1(n24020), .A2(n25653), .B1(n2121), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_5/N3 ) );
  AOI22_X1 U13107 ( .A1(n24011), .A2(n26772), .B1(n25148), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_11/N3 ) );
  AOI22_X1 U13058 ( .A1(n24010), .A2(n25609), .B1(n25156), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_11/N3 ) );
  AOI22_X1 U13277 ( .A1(n23996), .A2(n25652), .B1(n2118), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_5/N3 ) );
  AOI22_X1 U13320 ( .A1(n23996), .A2(n25604), .B1(n2694), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_1/N3 ) );
  AOI22_X1 U13009 ( .A1(n24010), .A2(n25655), .B1(n24953), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_6/N3 ) );
  AOI22_X1 U13216 ( .A1(n24020), .A2(n25605), .B1(n2697), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_1/N3 ) );
  AOI22_X1 U13150 ( .A1(n24001), .A2(n25622), .B1(n24939), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_19/N3 ) );
  AOI22_X1 U13201 ( .A1(n24020), .A2(n25623), .B1(n25133), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_19/N3 ) );
  AOI22_X1 U13164 ( .A1(n24001), .A2(n25604), .B1(n2696), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_1/N3 ) );
  AOI22_X1 U13073 ( .A1(n24011), .A2(n26748), .B1(n24673), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_6/N3 ) );
  AOI22_X1 U13459 ( .A1(n23998), .A2(n25656), .B1(n24778), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_7/N3 ) );
  AOI22_X1 U13438 ( .A1(n23999), .A2(n26769), .B1(n24898), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_15/N3 ) );
  AOI22_X1 U13319 ( .A1(n23996), .A2(n25606), .B1(n3054), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_10/N3 ) );
  AOI22_X1 U13330 ( .A1(n24000), .A2(n25655), .B1(n24593), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_6/N3 ) );
  AOI22_X1 U13396 ( .A1(n23999), .A2(n26748), .B1(n24917), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_6/N3 ) );
  AOI22_X1 U13215 ( .A1(n24020), .A2(n25607), .B1(n3057), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_10/N3 ) );
  AOI22_X1 U13120 ( .A1(n24001), .A2(n25656), .B1(n2048), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_7/N3 ) );
  AOI22_X1 U13171 ( .A1(n24020), .A2(n25657), .B1(n2049), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_7/N3 ) );
  AOI22_X1 U13296 ( .A1(n23996), .A2(n25630), .B1(n25070), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_23/N3 ) );
  AOI22_X1 U13071 ( .A1(n24011), .A2(n26747), .B1(n24662), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_7/N3 ) );
  AOI22_X1 U13163 ( .A1(n24001), .A2(n25606), .B1(n3056), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_10/N3 ) );
  AOI22_X1 U13109 ( .A1(n24011), .A2(n26773), .B1(n25147), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_10/N3 ) );
  AOI22_X1 U13461 ( .A1(n23998), .A2(n25654), .B1(n25106), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_6/N3 ) );
  AOI22_X1 U13007 ( .A1(n24010), .A2(n25657), .B1(n25042), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_7/N3 ) );
  AOI22_X1 U13005 ( .A1(n24010), .A2(n25659), .B1(n25043), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_8/N3 ) );
  AOI22_X1 U13394 ( .A1(n23999), .A2(n26747), .B1(n24918), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_7/N3 ) );
  AOI22_X1 U13064 ( .A1(n24010), .A2(n25603), .B1(n25153), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_0/N3 ) );
  AOI22_X1 U13478 ( .A1(n23998), .A2(n25627), .B1(n738), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_21/N3 ) );
  AOI22_X1 U13424 ( .A1(n23999), .A2(n26762), .B1(n24904), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_21/N3 ) );
  AOI22_X1 U13358 ( .A1(n24000), .A2(n25628), .B1(n25118), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_21/N3 ) );
  AOI22_X1 U13495 ( .A1(n23998), .A2(n25606), .B1(n25265), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_10/N3 ) );
  AOI22_X1 U13422 ( .A1(n23999), .A2(n26761), .B1(net741170), .B2(n20549), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_17/DFF_22/N3 ) );
  AOI22_X1 U13305 ( .A1(n23996), .A2(n25622), .B1(n25068), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_19/N3 ) );
  AOI22_X1 U13091 ( .A1(n24011), .A2(n26762), .B1(n741), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_21/N3 ) );
  AOI22_X1 U13113 ( .A1(n24011), .A2(n26775), .B1(n25145), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_0/N3 ) );
  AOI22_X1 U13497 ( .A1(n23998), .A2(n25604), .B1(n25264), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_1/N3 ) );
  AOI22_X1 U13036 ( .A1(n24010), .A2(n25628), .B1(n25164), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_21/N3 ) );
  AOI22_X1 U13450 ( .A1(n23999), .A2(n26774), .B1(n24893), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_1/N3 ) );
  AOI22_X1 U13386 ( .A1(n24000), .A2(n25603), .B1(n25107), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_0/N3 ) );
  AOI22_X1 U13384 ( .A1(n24000), .A2(n25605), .B1(n25108), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_1/N3 ) );
  AOI22_X1 U13034 ( .A1(n24010), .A2(n25629), .B1(net740886), .B2(n20400), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_23/DFF_22/N3 ) );
  AOI22_X1 U13111 ( .A1(n24011), .A2(n26774), .B1(n25146), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_1/N3 ) );
  AOI22_X1 U13448 ( .A1(n23999), .A2(n26773), .B1(n24894), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_10/N3 ) );
  AOI22_X1 U13090 ( .A1(n24011), .A2(n26761), .B1(n818), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_22/N3 ) );
  AOI22_X1 U13275 ( .A1(n23996), .A2(n25656), .B1(n2046), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_7/N3 ) );
  AOI22_X1 U13356 ( .A1(n24000), .A2(n25629), .B1(net740936), .B2(n20521), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_18/DFF_22/N3 ) );
  AOI22_X1 U13392 ( .A1(n23999), .A2(n26746), .B1(n24919), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_8/N3 ) );
  AOI22_X1 U13477 ( .A1(n23998), .A2(net717153), .B1(n815), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_22/N3 ) );
  AOI22_X1 U13062 ( .A1(n24010), .A2(n25605), .B1(n25154), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_1/N3 ) );
  AOI22_X1 U13382 ( .A1(n24000), .A2(n25607), .B1(n25109), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_10/N3 ) );
  AOI22_X1 U13452 ( .A1(n23999), .A2(n26775), .B1(n24892), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_0/N3 ) );
  AOI22_X1 U13089 ( .A1(n24011), .A2(n26760), .B1(n779), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_23/N3 ) );
  AOI22_X1 U13499 ( .A1(n23998), .A2(n25602), .B1(n25263), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_0/N3 ) );
  AOI22_X1 U13420 ( .A1(n23999), .A2(n26760), .B1(n24905), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_23/N3 ) );
  AOI22_X1 U13476 ( .A1(n23998), .A2(n25630), .B1(n776), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_23/N3 ) );
  AOI22_X1 U13192 ( .A1(n24020), .A2(n25631), .B1(n25135), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_23/N3 ) );
  AOI22_X1 U13060 ( .A1(n24010), .A2(n25607), .B1(n25155), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_10/N3 ) );
  AOI22_X1 U13141 ( .A1(n24001), .A2(n25630), .B1(n24941), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_23/N3 ) );
  AOI22_X1 U13069 ( .A1(n24011), .A2(n26746), .B1(n24666), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_8/N3 ) );
  AOI22_X1 U13326 ( .A1(n24000), .A2(n25659), .B1(n24590), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_8/N3 ) );
  AOI22_X1 U13298 ( .A1(n23996), .A2(net717153), .B1(net740989), .B2(n20502), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_19/DFF_22/N3 ) );
  AOI22_X1 U13170 ( .A1(n24020), .A2(n25659), .B1(n2013), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_8/N3 ) );
  AOI22_X1 U13119 ( .A1(n24001), .A2(n25658), .B1(n2012), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_8/N3 ) );
  AOI22_X1 U13321 ( .A1(n23996), .A2(n25602), .B1(n3090), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_0/N3 ) );
  AOI22_X1 U13143 ( .A1(n24001), .A2(net717153), .B1(net741130), .B2(n20445), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_21/DFF_22/N3 ) );
  AOI22_X1 U13274 ( .A1(n23996), .A2(n25658), .B1(n2010), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_8/N3 ) );
  AOI22_X1 U13276 ( .A1(n23996), .A2(n25654), .B1(n2082), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_6/N3 ) );
  AOI22_X1 U13172 ( .A1(n24020), .A2(n25655), .B1(n2085), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_6/N3 ) );
  AOI22_X1 U13217 ( .A1(n24020), .A2(n25603), .B1(n3098), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_0/N3 ) );
  AOI22_X1 U13194 ( .A1(n24020), .A2(n25629), .B1(net740918), .B2(n20464), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_20/DFF_22/N3 ) );
  AOI22_X1 U13165 ( .A1(n24001), .A2(n25602), .B1(n3097), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_0/N3 ) );
  AOI22_X1 U13457 ( .A1(n23998), .A2(n25658), .B1(n24779), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_8/N3 ) );
  AOI22_X1 U13121 ( .A1(n24001), .A2(n25654), .B1(n2084), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_6/N3 ) );
  AOI22_X1 U13354 ( .A1(n24000), .A2(n25631), .B1(n25119), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_23/N3 ) );
  AOI22_X1 U13032 ( .A1(n24010), .A2(n25631), .B1(n25165), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_23/N3 ) );
  AOI22_X1 U13052 ( .A1(n20398), .A2(n25613), .B1(n25158), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_14/N3 ) );
  AOI22_X1 U13338 ( .A1(n24000), .A2(n25647), .B1(n25126), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_30/N3 ) );
  AOI22_X1 U13159 ( .A1(n24001), .A2(n25612), .B1(n2912), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_14/N3 ) );
  AOI22_X1 U13016 ( .A1(n20398), .A2(n25647), .B1(n25172), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_30/N3 ) );
  AOI22_X1 U13126 ( .A1(n24001), .A2(n25646), .B1(n24948), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_30/N3 ) );
  AOI22_X1 U13210 ( .A1(n20462), .A2(n25613), .B1(n2913), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_14/N3 ) );
  AOI22_X1 U13314 ( .A1(n23996), .A2(n25612), .B1(n2910), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_14/N3 ) );
  AOI22_X1 U13487 ( .A1(n23998), .A2(n25612), .B1(n25267), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_14/N3 ) );
  AOI22_X1 U13101 ( .A1(n20432), .A2(n26770), .B1(n25150), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_14/N3 ) );
  AOI22_X1 U13374 ( .A1(n24000), .A2(n25613), .B1(n25112), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_14/N3 ) );
  AOI22_X1 U13080 ( .A1(n20432), .A2(n26752), .B1(n506), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_30/N3 ) );
  AOI22_X1 U13281 ( .A1(n23996), .A2(n25646), .B1(n25077), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_30/N3 ) );
  AOI22_X1 U13440 ( .A1(n23999), .A2(n26770), .B1(n24897), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_14/N3 ) );
  AOI22_X1 U13468 ( .A1(n23998), .A2(n25646), .B1(n503), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_30/N3 ) );
  AOI22_X1 U13404 ( .A1(n23999), .A2(n26752), .B1(n24913), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_30/N3 ) );
  AOI22_X1 U13177 ( .A1(n20462), .A2(n25647), .B1(n25142), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_30/N3 ) );
  AOI22_X1 U13129 ( .A1(n24001), .A2(n25642), .B1(n24947), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_29/N3 ) );
  AOI22_X1 U13180 ( .A1(n20462), .A2(n25643), .B1(n25141), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_29/N3 ) );
  AOI22_X1 U13288 ( .A1(n23996), .A2(n25638), .B1(n25074), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_27/N3 ) );
  AOI22_X1 U13184 ( .A1(n20462), .A2(n25639), .B1(n25139), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_27/N3 ) );
  AOI22_X1 U13133 ( .A1(n24001), .A2(n25638), .B1(n24945), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_27/N3 ) );
  AOI22_X1 U13020 ( .A1(n20398), .A2(n25643), .B1(n25171), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_29/N3 ) );
  AOI22_X1 U13083 ( .A1(n20432), .A2(n26754), .B1(n432), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_29/N3 ) );
  AOI22_X1 U13342 ( .A1(n24000), .A2(n25643), .B1(n25125), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_29/N3 ) );
  AOI22_X1 U13408 ( .A1(n23999), .A2(n26754), .B1(n24911), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_29/N3 ) );
  AOI22_X1 U13198 ( .A1(n20462), .A2(n25626), .B1(net740920), .B2(n20464), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_20/DFF_20/N3 ) );
  AOI22_X1 U13470 ( .A1(n23998), .A2(n25642), .B1(n429), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_29/N3 ) );
  AOI22_X1 U13147 ( .A1(n24001), .A2(net717157), .B1(net741132), .B2(n20445), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_21/DFF_20/N3 ) );
  AOI22_X1 U13472 ( .A1(n23998), .A2(n25638), .B1(n582), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_27/N3 ) );
  AOI22_X1 U13412 ( .A1(n23999), .A2(n26756), .B1(n24909), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_27/N3 ) );
  AOI22_X1 U13456 ( .A1(n23998), .A2(n25660), .B1(n353), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_9/N3 ) );
  AOI22_X1 U13346 ( .A1(n24000), .A2(n25639), .B1(n25123), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_27/N3 ) );
  AOI22_X1 U13085 ( .A1(n20432), .A2(n26756), .B1(n585), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_27/N3 ) );
  AOI22_X1 U13024 ( .A1(n20398), .A2(n25639), .B1(n25169), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_27/N3 ) );
  AOI22_X1 U13272 ( .A1(n23996), .A2(n25660), .B1(n24667), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_9/N3 ) );
  AOI22_X1 U13479 ( .A1(n23998), .A2(net717157), .B1(n855), .B2(n20582), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_20/N3 ) );
  AOI22_X1 U13426 ( .A1(n23999), .A2(n26763), .B1(net741172), .B2(n20549), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_17/DFF_20/N3 ) );
  AOI22_X1 U13168 ( .A1(n20462), .A2(n25661), .B1(n25144), .B2(n20464), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_9/N3 ) );
  AOI22_X1 U13117 ( .A1(n24001), .A2(n25660), .B1(n24950), .B2(n20445), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_9/N3 ) );
  AOI22_X1 U13284 ( .A1(n23996), .A2(n25642), .B1(n25076), .B2(n20502), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_29/N3 ) );
  AOI22_X1 U13360 ( .A1(n24000), .A2(n25626), .B1(net740938), .B2(n20521), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_18/DFF_20/N3 ) );
  AOI22_X1 U13092 ( .A1(n20432), .A2(n26763), .B1(n858), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_20/N3 ) );
  AOI22_X1 U13302 ( .A1(n23996), .A2(net717157), .B1(net740991), .B2(n20502), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_19/DFF_20/N3 ) );
  AOI22_X1 U13324 ( .A1(n24000), .A2(n25661), .B1(n25129), .B2(n20521), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_9/N3 ) );
  AOI22_X1 U13068 ( .A1(n20432), .A2(n26745), .B1(n356), .B2(n20433), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_9/N3 ) );
  AOI22_X1 U13003 ( .A1(n20398), .A2(n25661), .B1(n25173), .B2(n20400), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_9/N3 ) );
  AOI22_X1 U13038 ( .A1(n20398), .A2(n25626), .B1(net740888), .B2(n20400), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_23/DFF_20/N3 ) );
  AOI22_X1 U13390 ( .A1(n23999), .A2(n26745), .B1(n24920), .B2(n20549), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_9/N3 ) );
  AOI22_X1 U12224 ( .A1(n25673), .A2(n25653), .B1(n2140), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_5/N3 ) );
  AOI22_X1 U12231 ( .A1(n25673), .A2(n25643), .B1(n25032), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_29/N3 ) );
  AOI22_X1 U12219 ( .A1(n25673), .A2(n25661), .B1(n25035), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_9/N3 ) );
  AOI22_X1 U12239 ( .A1(n25673), .A2(n25635), .B1(n25028), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_25/N3 ) );
  AOI22_X1 U12223 ( .A1(n20134), .A2(n25655), .B1(n2104), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_6/N3 ) );
  AOI22_X1 U12264 ( .A1(n25673), .A2(n25609), .B1(n3040), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_11/N3 ) );
  AOI22_X1 U12221 ( .A1(n25673), .A2(n25659), .B1(n2032), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_8/N3 ) );
  AOI22_X1 U12261 ( .A1(n25673), .A2(n25613), .B1(n2932), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_14/N3 ) );
  AOI22_X1 U12265 ( .A1(n25673), .A2(n25607), .B1(n3076), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_10/N3 ) );
  AOI22_X1 U12225 ( .A1(n25673), .A2(n25651), .B1(n2176), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_4/N3 ) );
  AOI22_X1 U12226 ( .A1(n25673), .A2(n25649), .B1(n25034), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_31/N3 ) );
  AOI22_X1 U12245 ( .A1(n25673), .A2(n25629), .B1(net741037), .B2(n25672), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_9/DFF_22/N3 ) );
  AOI22_X1 U12267 ( .A1(n20134), .A2(n25603), .B1(n3131), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_0/N3 ) );
  AOI22_X1 U12256 ( .A1(n25673), .A2(n25619), .B1(n25022), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_17/N3 ) );
  AOI22_X1 U12266 ( .A1(n25673), .A2(n25605), .B1(n2716), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_1/N3 ) );
  AOI22_X1 U12228 ( .A1(n25673), .A2(n25647), .B1(n25033), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_30/N3 ) );
  AOI22_X1 U12260 ( .A1(n25673), .A2(n25615), .B1(n2896), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_15/N3 ) );
  AOI22_X1 U12254 ( .A1(n25673), .A2(n25621), .B1(n25023), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_18/N3 ) );
  AOI22_X1 U12251 ( .A1(n25673), .A2(n25625), .B1(n2320), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_2/N3 ) );
  AOI22_X1 U12237 ( .A1(n25673), .A2(n25637), .B1(n25029), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_26/N3 ) );
  AOI22_X1 U12230 ( .A1(n25673), .A2(n25645), .B1(n2212), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_3/N3 ) );
  AOI22_X1 U12235 ( .A1(n25673), .A2(n25639), .B1(n25030), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_27/N3 ) );
  AOI22_X1 U12243 ( .A1(n25673), .A2(n25631), .B1(n25026), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_23/N3 ) );
  AOI22_X1 U12249 ( .A1(n25673), .A2(n25626), .B1(net741039), .B2(n25672), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_9/DFF_20/N3 ) );
  AOI22_X1 U12241 ( .A1(n25673), .A2(n25633), .B1(n25027), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_24/N3 ) );
  AOI22_X1 U12222 ( .A1(n25673), .A2(n25657), .B1(n2068), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_7/N3 ) );
  AOI22_X1 U12262 ( .A1(n25673), .A2(n25611), .B1(n2968), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_13/N3 ) );
  AOI22_X1 U12252 ( .A1(n25673), .A2(n25623), .B1(n25024), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_19/N3 ) );
  AOI22_X1 U12258 ( .A1(n25673), .A2(n25617), .B1(n25021), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_16/N3 ) );
  AOI22_X1 U12247 ( .A1(n25673), .A2(n25628), .B1(n25025), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_21/N3 ) );
  AOI22_X1 U12233 ( .A1(n20134), .A2(n25641), .B1(n25031), .B2(n25672), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_28/N3 ) );
  AOI22_X1 U12328 ( .A1(n25671), .A2(n26773), .B1(n25001), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_10/N3 ) );
  AOI22_X1 U12307 ( .A1(n25671), .A2(n26764), .B1(n24674), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_2/N3 ) );
  AOI22_X1 U12326 ( .A1(n25671), .A2(n26772), .B1(n25002), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_11/N3 ) );
  AOI22_X1 U12330 ( .A1(n25671), .A2(n26774), .B1(n25000), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_1/N3 ) );
  AOI22_X1 U12332 ( .A1(n20155), .A2(n26775), .B1(n24999), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_0/N3 ) );
  AOI22_X1 U12301 ( .A1(n25671), .A2(n26761), .B1(net741054), .B2(n25670), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_8/DFF_22/N3 ) );
  AOI22_X1 U12291 ( .A1(n25671), .A2(n26756), .B1(n25015), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_27/N3 ) );
  AOI22_X1 U12311 ( .A1(n25671), .A2(n26766), .B1(n25008), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_18/N3 ) );
  AOI22_X1 U12295 ( .A1(n25671), .A2(n26758), .B1(n25013), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_25/N3 ) );
  AOI22_X1 U12299 ( .A1(n25671), .A2(n26760), .B1(n25011), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_23/N3 ) );
  AOI22_X1 U12272 ( .A1(n25671), .A2(n26746), .B1(n24663), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_8/N3 ) );
  AOI22_X1 U12313 ( .A1(n25671), .A2(n26767), .B1(n25007), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_17/N3 ) );
  AOI22_X1 U12270 ( .A1(n25671), .A2(n26745), .B1(n25020), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_9/N3 ) );
  AOI22_X1 U12293 ( .A1(n25671), .A2(n26757), .B1(n25014), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_26/N3 ) );
  AOI22_X1 U12276 ( .A1(n25671), .A2(n26748), .B1(n24671), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_6/N3 ) );
  AOI22_X1 U12303 ( .A1(n25671), .A2(n26762), .B1(n25010), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_21/N3 ) );
  AOI22_X1 U12297 ( .A1(n25671), .A2(n26759), .B1(n25012), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_24/N3 ) );
  AOI22_X1 U12287 ( .A1(n25671), .A2(n26754), .B1(n25017), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_29/N3 ) );
  AOI22_X1 U12309 ( .A1(n20155), .A2(n26765), .B1(n25009), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_19/N3 ) );
  AOI22_X1 U12278 ( .A1(n25671), .A2(n26749), .B1(n24668), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_5/N3 ) );
  AOI22_X1 U12305 ( .A1(n20155), .A2(n26763), .B1(net741056), .B2(n25670), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_8/DFF_20/N3 ) );
  AOI22_X1 U12274 ( .A1(n25671), .A2(n26747), .B1(n24659), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_7/N3 ) );
  AOI22_X1 U12316 ( .A1(n25671), .A2(n26768), .B1(n25006), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_16/N3 ) );
  AOI22_X1 U12322 ( .A1(n25671), .A2(n26771), .B1(n25003), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_13/N3 ) );
  AOI22_X1 U12285 ( .A1(n25671), .A2(n26753), .B1(n24649), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_3/N3 ) );
  AOI22_X1 U12283 ( .A1(n25671), .A2(n26752), .B1(n25018), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_30/N3 ) );
  AOI22_X1 U12318 ( .A1(n25671), .A2(n26769), .B1(n25005), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_15/N3 ) );
  AOI22_X1 U12320 ( .A1(n25671), .A2(n26770), .B1(n25004), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_14/N3 ) );
  AOI22_X1 U12280 ( .A1(n25671), .A2(n26750), .B1(n25019), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_4/N3 ) );
  AOI22_X1 U12289 ( .A1(n25671), .A2(n26755), .B1(n25016), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_28/N3 ) );
  AOI22_X1 U12282 ( .A1(n25671), .A2(n26751), .B1(n475), .B2(n25670), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_31/N3 ) );
  AOI22_X1 U12533 ( .A1(n24017), .A2(n25606), .B1(n3069), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_10/N3 ) );
  AOI22_X1 U12513 ( .A1(n24017), .A2(net717153), .B1(net740818), .B2(n20243), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_4/DFF_22/N3 ) );
  AOI22_X1 U12520 ( .A1(n24017), .A2(n25622), .B1(n25225), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_19/N3 ) );
  AOI22_X1 U12535 ( .A1(n24017), .A2(n25602), .B1(n3117), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_0/N3 ) );
  AOI22_X1 U12509 ( .A1(n24017), .A2(n25632), .B1(n25228), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_24/N3 ) );
  AOI22_X1 U12501 ( .A1(n24017), .A2(n25640), .B1(n25232), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_28/N3 ) );
  AOI22_X1 U12528 ( .A1(n24017), .A2(n25614), .B1(n2889), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_15/N3 ) );
  AOI22_X1 U12534 ( .A1(n24017), .A2(n25604), .B1(n2709), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_1/N3 ) );
  AOI22_X1 U12524 ( .A1(n24017), .A2(n25618), .B1(n25223), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_17/N3 ) );
  AOI22_X1 U12498 ( .A1(n24017), .A2(n25644), .B1(n2205), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_3/N3 ) );
  AOI22_X1 U12511 ( .A1(n24017), .A2(n25630), .B1(n25227), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_23/N3 ) );
  AOI22_X1 U12493 ( .A1(n24017), .A2(n25650), .B1(n2169), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_4/N3 ) );
  AOI22_X1 U12490 ( .A1(n24017), .A2(n25656), .B1(n2061), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_7/N3 ) );
  AOI22_X1 U12505 ( .A1(n24017), .A2(n25636), .B1(n25230), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_26/N3 ) );
  AOI22_X1 U12507 ( .A1(n24017), .A2(n25634), .B1(n25229), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_25/N3 ) );
  AOI22_X1 U12491 ( .A1(n24017), .A2(n25654), .B1(n2097), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_6/N3 ) );
  AOI22_X1 U12532 ( .A1(n24017), .A2(n25608), .B1(n3033), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_11/N3 ) );
  AOI22_X1 U12522 ( .A1(n24017), .A2(n25620), .B1(n25224), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_18/N3 ) );
  AOI22_X1 U12489 ( .A1(n24017), .A2(n25658), .B1(n2025), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_8/N3 ) );
  AOI22_X1 U12526 ( .A1(n24017), .A2(n25616), .B1(n25222), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_16/N3 ) );
  AOI22_X1 U12530 ( .A1(n24017), .A2(n25610), .B1(n2961), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_13/N3 ) );
  AOI22_X1 U12494 ( .A1(n24017), .A2(n25648), .B1(n25235), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_31/N3 ) );
  AOI22_X1 U12519 ( .A1(n24017), .A2(n25624), .B1(n2313), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_2/N3 ) );
  AOI22_X1 U12492 ( .A1(n24017), .A2(n25652), .B1(n2133), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_5/N3 ) );
  AOI22_X1 U12515 ( .A1(n24017), .A2(n25627), .B1(n25226), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_21/N3 ) );
  AOI22_X1 U12468 ( .A1(n24016), .A2(n26764), .B1(n2317), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_2/N3 ) );
  AOI22_X1 U12469 ( .A1(n24016), .A2(n26765), .B1(n25053), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_19/N3 ) );
  AOI22_X1 U12477 ( .A1(n24016), .A2(n26769), .B1(n2893), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_15/N3 ) );
  AOI22_X1 U12440 ( .A1(n24016), .A2(n26748), .B1(n2101), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_6/N3 ) );
  AOI22_X1 U12450 ( .A1(n24016), .A2(n26755), .B1(n25060), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_28/N3 ) );
  AOI22_X1 U12441 ( .A1(n24016), .A2(n26749), .B1(n2137), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_5/N3 ) );
  AOI22_X1 U12481 ( .A1(n24016), .A2(n26772), .B1(n3037), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_11/N3 ) );
  AOI22_X1 U12471 ( .A1(n24016), .A2(n26766), .B1(n25052), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_18/N3 ) );
  AOI22_X1 U12473 ( .A1(n24016), .A2(n26767), .B1(n25051), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_17/N3 ) );
  AOI22_X1 U12464 ( .A1(n24016), .A2(n26762), .B1(n25054), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_21/N3 ) );
  AOI22_X1 U12442 ( .A1(n24016), .A2(n26750), .B1(n2173), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_4/N3 ) );
  AOI22_X1 U12438 ( .A1(n24016), .A2(n26746), .B1(n2029), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_8/N3 ) );
  AOI22_X1 U12462 ( .A1(n24016), .A2(n26761), .B1(net741006), .B2(n20223), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_5/DFF_22/N3 ) );
  AOI22_X1 U12454 ( .A1(n24016), .A2(n26757), .B1(n25058), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_26/N3 ) );
  AOI22_X1 U12482 ( .A1(n24016), .A2(n26773), .B1(n3073), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_10/N3 ) );
  AOI22_X1 U12456 ( .A1(n24016), .A2(n26758), .B1(n25057), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_25/N3 ) );
  AOI22_X1 U12447 ( .A1(n24016), .A2(n26753), .B1(n2209), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_3/N3 ) );
  AOI22_X1 U12483 ( .A1(n24016), .A2(n26774), .B1(n2713), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_1/N3 ) );
  AOI22_X1 U12439 ( .A1(n24016), .A2(n26747), .B1(n2065), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_7/N3 ) );
  AOI22_X1 U12475 ( .A1(n24016), .A2(n26768), .B1(n25050), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_16/N3 ) );
  AOI22_X1 U12458 ( .A1(n24016), .A2(n26759), .B1(n25056), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_24/N3 ) );
  AOI22_X1 U12484 ( .A1(n24016), .A2(n26775), .B1(n3125), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_0/N3 ) );
  AOI22_X1 U12460 ( .A1(n24016), .A2(n26760), .B1(n25055), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_23/N3 ) );
  AOI22_X1 U12479 ( .A1(n24016), .A2(n26771), .B1(n2965), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_13/N3 ) );
  AOI22_X1 U12443 ( .A1(n24016), .A2(n26751), .B1(n25063), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_31/N3 ) );
  AOI22_X1 U12430 ( .A1(n24015), .A2(n25609), .B1(n3036), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_11/N3 ) );
  AOI22_X1 U12433 ( .A1(n24015), .A2(n25603), .B1(n3124), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_0/N3 ) );
  AOI22_X1 U12405 ( .A1(n24015), .A2(n25635), .B1(n25244), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_25/N3 ) );
  AOI22_X1 U12407 ( .A1(n24015), .A2(n25633), .B1(n25243), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_24/N3 ) );
  AOI22_X1 U12428 ( .A1(n24015), .A2(n25611), .B1(n2964), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_13/N3 ) );
  AOI22_X1 U12409 ( .A1(n24015), .A2(n25631), .B1(n25242), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_23/N3 ) );
  AOI22_X1 U12403 ( .A1(n24015), .A2(n25637), .B1(n25245), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_26/N3 ) );
  AOI22_X1 U12389 ( .A1(n24015), .A2(n25655), .B1(n2100), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_6/N3 ) );
  AOI22_X1 U12426 ( .A1(n24015), .A2(n25615), .B1(n2892), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_15/N3 ) );
  AOI22_X1 U12390 ( .A1(n24015), .A2(n25653), .B1(n2136), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_5/N3 ) );
  AOI22_X1 U12418 ( .A1(n24015), .A2(n25623), .B1(n25240), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_19/N3 ) );
  AOI22_X1 U12399 ( .A1(n24015), .A2(n25641), .B1(n25247), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_28/N3 ) );
  AOI22_X1 U12391 ( .A1(n24015), .A2(n25651), .B1(n2172), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_4/N3 ) );
  AOI22_X1 U12411 ( .A1(n24015), .A2(n25629), .B1(net740801), .B2(n20204), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_6/DFF_22/N3 ) );
  AOI22_X1 U12387 ( .A1(n24015), .A2(n25659), .B1(n2028), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_8/N3 ) );
  AOI22_X1 U12396 ( .A1(n24015), .A2(n25645), .B1(n2208), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_3/N3 ) );
  AOI22_X1 U12392 ( .A1(n24015), .A2(n25649), .B1(n24656), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_31/N3 ) );
  AOI22_X1 U12413 ( .A1(n24015), .A2(n25628), .B1(n25241), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_21/N3 ) );
  AOI22_X1 U12431 ( .A1(n24015), .A2(n25607), .B1(n3072), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_10/N3 ) );
  AOI22_X1 U12422 ( .A1(n24015), .A2(n25619), .B1(n25238), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_17/N3 ) );
  AOI22_X1 U12388 ( .A1(n24015), .A2(n25657), .B1(n2064), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_7/N3 ) );
  AOI22_X1 U12432 ( .A1(n24015), .A2(n25605), .B1(n2712), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_1/N3 ) );
  AOI22_X1 U12420 ( .A1(n24015), .A2(n25621), .B1(n25239), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_18/N3 ) );
  AOI22_X1 U12417 ( .A1(n24015), .A2(n25625), .B1(n2316), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_2/N3 ) );
  AOI22_X1 U12424 ( .A1(n24015), .A2(n25617), .B1(n25237), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_16/N3 ) );
  AOI22_X1 U12496 ( .A1(n20241), .A2(n25646), .B1(n25234), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_30/N3 ) );
  AOI22_X1 U12517 ( .A1(n20241), .A2(net717157), .B1(net740820), .B2(n20243), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_4/DFF_20/N3 ) );
  AOI22_X1 U12487 ( .A1(n20241), .A2(n25660), .B1(n25236), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_9/N3 ) );
  AOI22_X1 U12529 ( .A1(n20241), .A2(n25612), .B1(n2925), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_14/N3 ) );
  AOI22_X1 U12503 ( .A1(n20241), .A2(n25638), .B1(n25231), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_27/N3 ) );
  AOI22_X1 U12499 ( .A1(n20241), .A2(n25642), .B1(n25233), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_29/N3 ) );
  AOI22_X1 U12436 ( .A1(n20221), .A2(n26745), .B1(n25064), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_9/N3 ) );
  AOI22_X1 U12478 ( .A1(n20221), .A2(n26770), .B1(n2929), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_14/N3 ) );
  AOI22_X1 U12448 ( .A1(n20221), .A2(n26754), .B1(n25061), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_29/N3 ) );
  AOI22_X1 U12445 ( .A1(n20221), .A2(n26752), .B1(n25062), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_30/N3 ) );
  AOI22_X1 U12466 ( .A1(n20221), .A2(n26763), .B1(net741008), .B2(n20223), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_5/DFF_20/N3 ) );
  AOI22_X1 U12452 ( .A1(n20221), .A2(n26756), .B1(n25059), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_27/N3 ) );
  AOI22_X1 U12394 ( .A1(n20202), .A2(n25647), .B1(n25249), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_30/N3 ) );
  AOI22_X1 U12415 ( .A1(n20202), .A2(n25626), .B1(net740803), .B2(n20204), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_6/DFF_20/N3 ) );
  AOI22_X1 U12397 ( .A1(n20202), .A2(n25643), .B1(n25248), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_29/N3 ) );
  AOI22_X1 U12401 ( .A1(n20202), .A2(n25639), .B1(n25246), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_27/N3 ) );
  AOI22_X1 U12385 ( .A1(n20202), .A2(n25661), .B1(n25079), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_9/N3 ) );
  AOI22_X1 U12427 ( .A1(n20202), .A2(n25613), .B1(n2928), .B2(n20204), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_14/N3 ) );
  AOI22_X1 U12686 ( .A1(n24019), .A2(n25624), .B1(n2314), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_2/N3 ) );
  AOI22_X1 U12702 ( .A1(n24019), .A2(n25602), .B1(n3118), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_0/N3 ) );
  AOI22_X1 U12659 ( .A1(n24019), .A2(n25652), .B1(n2134), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_5/N3 ) );
  AOI22_X1 U12701 ( .A1(n24019), .A2(n25604), .B1(n2710), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_1/N3 ) );
  AOI22_X1 U12660 ( .A1(n24019), .A2(n25650), .B1(n2170), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_4/N3 ) );
  AOI22_X1 U12665 ( .A1(n24019), .A2(n25644), .B1(n2206), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_3/N3 ) );
  AOI22_X1 U12658 ( .A1(n24019), .A2(n25654), .B1(n2098), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_6/N3 ) );
  AOI22_X1 U12676 ( .A1(n24019), .A2(n25632), .B1(n24990), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_24/N3 ) );
  AOI22_X1 U12687 ( .A1(n24019), .A2(n25622), .B1(n24987), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_19/N3 ) );
  AOI22_X1 U12661 ( .A1(n24019), .A2(n25648), .B1(n24997), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_31/N3 ) );
  AOI22_X1 U12680 ( .A1(n24019), .A2(net717153), .B1(net741078), .B2(n20315), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_3/DFF_22/N3 ) );
  AOI22_X1 U12682 ( .A1(n24019), .A2(n25627), .B1(n24988), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_21/N3 ) );
  AOI22_X1 U12678 ( .A1(n24019), .A2(n25630), .B1(n24989), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_23/N3 ) );
  AOI22_X1 U12668 ( .A1(n24019), .A2(n25640), .B1(n24994), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_28/N3 ) );
  AOI22_X1 U12656 ( .A1(n24019), .A2(n25658), .B1(n2026), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_8/N3 ) );
  AOI22_X1 U12672 ( .A1(n24019), .A2(n25636), .B1(n24992), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_26/N3 ) );
  AOI22_X1 U12700 ( .A1(n24019), .A2(n25606), .B1(n3070), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_10/N3 ) );
  AOI22_X1 U12699 ( .A1(n24019), .A2(n25608), .B1(n3034), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_11/N3 ) );
  AOI22_X1 U12697 ( .A1(n24019), .A2(n25610), .B1(n2962), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_13/N3 ) );
  AOI22_X1 U12674 ( .A1(n24019), .A2(n25634), .B1(n24991), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_25/N3 ) );
  AOI22_X1 U12689 ( .A1(n24019), .A2(n25620), .B1(n24986), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_18/N3 ) );
  AOI22_X1 U12693 ( .A1(n24019), .A2(n25616), .B1(n24984), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_16/N3 ) );
  AOI22_X1 U12695 ( .A1(n24019), .A2(n25614), .B1(n2890), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_15/N3 ) );
  AOI22_X1 U12691 ( .A1(n24019), .A2(n25618), .B1(n24985), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_17/N3 ) );
  AOI22_X1 U12657 ( .A1(n24019), .A2(n25656), .B1(n2062), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_7/N3 ) );
  AOI22_X1 U13227 ( .A1(n24021), .A2(n26751), .B1(n24934), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_31/N3 ) );
  AOI22_X1 U13252 ( .A1(n24021), .A2(n26764), .B1(n2307), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_2/N3 ) );
  AOI22_X1 U13246 ( .A1(n24021), .A2(n26761), .B1(net741147), .B2(n20483), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_2/DFF_22/N3 ) );
  AOI22_X1 U13269 ( .A1(n24021), .A2(n26775), .B1(n3108), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_0/N3 ) );
  AOI22_X1 U13248 ( .A1(n24021), .A2(n26762), .B1(n24925), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_21/N3 ) );
  AOI22_X1 U13242 ( .A1(n24021), .A2(n26759), .B1(n24927), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_24/N3 ) );
  AOI22_X1 U13234 ( .A1(n24021), .A2(n26755), .B1(n24931), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_28/N3 ) );
  AOI22_X1 U13253 ( .A1(n24021), .A2(n26765), .B1(n24924), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_19/N3 ) );
  AOI22_X1 U13267 ( .A1(n24021), .A2(n26773), .B1(n3063), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_10/N3 ) );
  AOI22_X1 U13224 ( .A1(n24021), .A2(n26748), .B1(n2091), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_6/N3 ) );
  AOI22_X1 U13259 ( .A1(n24021), .A2(n26768), .B1(n24921), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_16/N3 ) );
  AOI22_X1 U13244 ( .A1(n24021), .A2(n26760), .B1(n24926), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_23/N3 ) );
  AOI22_X1 U13261 ( .A1(n24021), .A2(n26769), .B1(n2883), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_15/N3 ) );
  AOI22_X1 U13263 ( .A1(n24021), .A2(n26771), .B1(n25078), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_13/N3 ) );
  AOI22_X1 U13222 ( .A1(n24021), .A2(n26746), .B1(n2019), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_8/N3 ) );
  AOI22_X1 U13231 ( .A1(n24021), .A2(n26753), .B1(n2199), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_3/N3 ) );
  AOI22_X1 U13226 ( .A1(n24021), .A2(n26750), .B1(n2163), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_4/N3 ) );
  AOI22_X1 U13238 ( .A1(n24021), .A2(n26757), .B1(n24929), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_26/N3 ) );
  AOI22_X1 U13257 ( .A1(n24021), .A2(n26767), .B1(n24922), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_17/N3 ) );
  AOI22_X1 U13268 ( .A1(n24021), .A2(n26774), .B1(n2703), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_1/N3 ) );
  AOI22_X1 U13240 ( .A1(n24021), .A2(n26758), .B1(n24928), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_25/N3 ) );
  AOI22_X1 U13255 ( .A1(n24021), .A2(n26766), .B1(n24923), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_18/N3 ) );
  AOI22_X1 U13225 ( .A1(n24021), .A2(n26749), .B1(n2127), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_5/N3 ) );
  AOI22_X1 U13266 ( .A1(n24021), .A2(n26772), .B1(n3027), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_11/N3 ) );
  AOI22_X1 U13223 ( .A1(n24021), .A2(n26747), .B1(n2055), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_7/N3 ) );
  AOI22_X1 U12684 ( .A1(n20313), .A2(net717157), .B1(net741080), .B2(n20315), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_3/DFF_20/N3 ) );
  AOI22_X1 U12654 ( .A1(n20313), .A2(n25660), .B1(n24998), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_9/N3 ) );
  AOI22_X1 U12670 ( .A1(n20313), .A2(n25638), .B1(n24993), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_27/N3 ) );
  AOI22_X1 U12666 ( .A1(n20313), .A2(n25642), .B1(n24995), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_29/N3 ) );
  AOI22_X1 U12663 ( .A1(n20313), .A2(n25646), .B1(n24996), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_30/N3 ) );
  AOI22_X1 U12696 ( .A1(n20313), .A2(n25612), .B1(n2926), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_14/N3 ) );
  AOI22_X1 U13250 ( .A1(n20481), .A2(n26763), .B1(net741149), .B2(n20483), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_2/DFF_20/N3 ) );
  AOI22_X1 U13220 ( .A1(n20481), .A2(n26745), .B1(n24935), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_9/N3 ) );
  AOI22_X1 U13236 ( .A1(n20481), .A2(n26756), .B1(n24930), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_27/N3 ) );
  AOI22_X1 U13232 ( .A1(n20481), .A2(n26754), .B1(n24932), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_29/N3 ) );
  AOI22_X1 U13229 ( .A1(n20481), .A2(n26752), .B1(n24933), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_30/N3 ) );
  AOI22_X1 U13262 ( .A1(n20481), .A2(n26770), .B1(n2919), .B2(n20483), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_14/N3 ) );
  AOI22_X1 U13881 ( .A1(n24023), .A2(n25625), .B1(n2297), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_2/N3 ) );
  AOI22_X1 U13927 ( .A1(n24023), .A2(n25603), .B1(n3089), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_0/N3 ) );
  AOI22_X1 U13865 ( .A1(n24023), .A2(n25631), .B1(n25295), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_23/N3 ) );
  AOI22_X1 U13920 ( .A1(n24023), .A2(n25607), .B1(n3053), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_10/N3 ) );
  AOI22_X1 U13853 ( .A1(n24023), .A2(n25637), .B1(n25298), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_26/N3 ) );
  AOI22_X1 U13869 ( .A1(n24023), .A2(n25629), .B1(net740739), .B2(n20706), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_1/DFF_22/N3 ) );
  AOI22_X1 U13893 ( .A1(n24023), .A2(n25619), .B1(n25291), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_17/N3 ) );
  AOI22_X1 U13917 ( .A1(n24023), .A2(n25609), .B1(n3017), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_11/N3 ) );
  AOI22_X1 U13903 ( .A1(n24023), .A2(n25615), .B1(n2873), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_15/N3 ) );
  AOI22_X1 U13884 ( .A1(n24023), .A2(n25623), .B1(n25293), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_19/N3 ) );
  AOI22_X1 U13861 ( .A1(n24023), .A2(n25633), .B1(n25296), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_24/N3 ) );
  AOI22_X1 U13857 ( .A1(n24023), .A2(n25635), .B1(n25297), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_25/N3 ) );
  AOI22_X1 U13825 ( .A1(n24023), .A2(n25651), .B1(n2153), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_4/N3 ) );
  AOI22_X1 U13889 ( .A1(n24023), .A2(n25621), .B1(n25292), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_18/N3 ) );
  AOI22_X1 U13823 ( .A1(n24023), .A2(n25653), .B1(n2117), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_5/N3 ) );
  AOI22_X1 U13843 ( .A1(n24023), .A2(n25641), .B1(n25300), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_28/N3 ) );
  AOI22_X1 U13815 ( .A1(n24023), .A2(n25659), .B1(n2009), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_8/N3 ) );
  AOI22_X1 U13873 ( .A1(n24023), .A2(n25628), .B1(n25294), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_21/N3 ) );
  AOI22_X1 U13828 ( .A1(n24023), .A2(n25649), .B1(n24848), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_31/N3 ) );
  AOI22_X1 U13898 ( .A1(n24023), .A2(n25617), .B1(n25290), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_16/N3 ) );
  AOI22_X1 U13909 ( .A1(n24023), .A2(n25611), .B1(n24847), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_13/N3 ) );
  AOI22_X1 U13818 ( .A1(n24023), .A2(n25657), .B1(n2045), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_7/N3 ) );
  AOI22_X1 U13836 ( .A1(n24023), .A2(n25645), .B1(n2189), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_3/N3 ) );
  AOI22_X1 U13820 ( .A1(n24023), .A2(n25655), .B1(n2081), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_6/N3 ) );
  AOI22_X1 U13923 ( .A1(n24023), .A2(n25605), .B1(n2693), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_1/N3 ) );
  AOI22_X1 U13906 ( .A1(n20704), .A2(n25613), .B1(n2909), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_14/N3 ) );
  AOI22_X1 U13832 ( .A1(n20704), .A2(n25647), .B1(n25302), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_30/N3 ) );
  AOI22_X1 U13877 ( .A1(n20704), .A2(n25626), .B1(net740741), .B2(n20706), 
        .ZN(\core_inst/ID/REGISTER_FILE/REG_1/DFF_20/N3 ) );
  AOI22_X1 U13848 ( .A1(n20704), .A2(n25639), .B1(n25299), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_27/N3 ) );
  AOI22_X1 U13811 ( .A1(n20704), .A2(n25661), .B1(n24849), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_9/N3 ) );
  AOI22_X1 U13839 ( .A1(n20704), .A2(n25643), .B1(n25301), .B2(n20706), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_29/N3 ) );
  AOI22_X1 U12379 ( .A1(n25669), .A2(n25604), .B1(n25251), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_1/N3 ) );
  AOI22_X1 U12356 ( .A1(n25669), .A2(n25632), .B1(n671), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_24/N3 ) );
  AOI22_X1 U12381 ( .A1(n20183), .A2(n25602), .B1(n25250), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_0/N3 ) );
  AOI22_X1 U12365 ( .A1(n25669), .A2(n25618), .B1(n710), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_17/N3 ) );
  AOI22_X1 U12358 ( .A1(n25669), .A2(net717153), .B1(n825), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_22/N3 ) );
  AOI22_X1 U12359 ( .A1(n25669), .A2(n25627), .B1(n748), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_21/N3 ) );
  AOI22_X1 U12360 ( .A1(n25669), .A2(net717157), .B1(n865), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_20/N3 ) );
  AOI22_X1 U12357 ( .A1(n25669), .A2(n25630), .B1(n786), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_23/N3 ) );
  AOI22_X1 U12375 ( .A1(n25669), .A2(n25608), .B1(n25253), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_11/N3 ) );
  AOI22_X1 U12339 ( .A1(n25669), .A2(n25656), .B1(n25258), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_7/N3 ) );
  AOI22_X1 U12363 ( .A1(n25669), .A2(n25622), .B1(n904), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_19/N3 ) );
  AOI22_X1 U12361 ( .A1(n25669), .A2(n25624), .B1(n25314), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_2/N3 ) );
  AOI22_X1 U12353 ( .A1(n20183), .A2(n25638), .B1(n592), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_27/N3 ) );
  AOI22_X1 U12364 ( .A1(n25669), .A2(n25620), .B1(n943), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_18/N3 ) );
  AOI22_X1 U12352 ( .A1(n25669), .A2(n25640), .B1(n553), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_28/N3 ) );
  AOI22_X1 U12349 ( .A1(n25669), .A2(n25644), .B1(n25257), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_3/N3 ) );
  AOI22_X1 U12366 ( .A1(n25669), .A2(n25616), .B1(n983), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_16/N3 ) );
  AOI22_X1 U12367 ( .A1(n25669), .A2(n25614), .B1(n25256), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_15/N3 ) );
  AOI22_X1 U12371 ( .A1(n25669), .A2(n25610), .B1(n25254), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_13/N3 ) );
  AOI22_X1 U12336 ( .A1(n25669), .A2(n25660), .B1(n363), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_9/N3 ) );
  AOI22_X1 U12348 ( .A1(n25669), .A2(n25646), .B1(n513), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_30/N3 ) );
  AOI22_X1 U12345 ( .A1(n25669), .A2(n25650), .B1(n25045), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_4/N3 ) );
  AOI22_X1 U12343 ( .A1(n25669), .A2(n25652), .B1(n25288), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_5/N3 ) );
  AOI22_X1 U12351 ( .A1(n25669), .A2(n25642), .B1(n439), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_29/N3 ) );
  AOI22_X1 U12355 ( .A1(n25669), .A2(n25634), .B1(n401), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_25/N3 ) );
  AOI22_X1 U12347 ( .A1(n25669), .A2(n25648), .B1(n474), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_31/N3 ) );
  AOI22_X1 U12369 ( .A1(n25669), .A2(n25612), .B1(n25255), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_14/N3 ) );
  AOI22_X1 U12341 ( .A1(n20183), .A2(n25654), .B1(n25289), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_6/N3 ) );
  AOI22_X1 U12337 ( .A1(n25669), .A2(n25658), .B1(n25259), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_8/N3 ) );
  AOI22_X1 U12377 ( .A1(n25669), .A2(n25606), .B1(n25252), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_10/N3 ) );
  AOI22_X1 U12354 ( .A1(n25669), .A2(n25636), .B1(n631), .B2(n25668), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_26/N3 ) );
  NOR2_X1 U10131 ( .A1(n24680), .A2(n18139), .ZN(n18156) );
  NAND2_X1 U10136 ( .A1(s_IFID_IR[30]), .A2(n24813), .ZN(n18159) );
  NOR2_X1 U10135 ( .A1(n18187), .A2(n18188), .ZN(n18162) );
  OAI21_X1 U10111 ( .B1(n24584), .B2(n18132), .A(n18135), .ZN(
        \cu_inst/EX/DFF_4/N3 ) );
  OAI21_X1 U10109 ( .B1(s_IFID_IR[28]), .B2(n18132), .A(n18133), .ZN(
        \cu_inst/EX/DFF_6/N3 ) );
  OAI21_X1 U10107 ( .B1(s_IFID_IR[30]), .B2(n26779), .A(n18129), .ZN(
        \cu_inst/EX/DFF_9/N3 ) );
  NOR2_X1 U10110 ( .A1(s_IFID_IR[26]), .A2(n18132), .ZN(\cu_inst/EX/DFF_5/N3 )
         );
  NOR2_X1 U10113 ( .A1(n18138), .A2(n26779), .ZN(\cu_inst/EX/DFF_18/N3 ) );
  NAND2_X1 U10206 ( .A1(s_MEM_LOAD_TYPE[1]), .A2(s_MEM_LOAD_TYPE[0]), .ZN(
        n18200) );
  NOR2_X2 U12018 ( .A1(n20070), .A2(n20068), .ZN(n19335) );
  NAND3_X1 U15895 ( .A1(n19289), .A2(n19294), .A3(n19292), .ZN(n20182) );
  NOR2_X2 U10187 ( .A1(s_MEM_LOAD_TYPE[1]), .A2(s_MEM_LOAD_TYPE[0]), .ZN(
        n18203) );
  NAND2_X1 U11122 ( .A1(n19240), .A2(n19256), .ZN(n18387) );
  NOR2_X1 U11096 ( .A1(n19248), .A2(n19243), .ZN(n18325) );
  NOR2_X1 U12011 ( .A1(n20069), .A2(n20065), .ZN(n19332) );
  NOR2_X1 U11130 ( .A1(s_IFID_IR[16]), .A2(s_IFID_IR[20]), .ZN(n19239) );
  NAND2_X1 U11126 ( .A1(s_IFID_IR[16]), .A2(net741525), .ZN(n19248) );
  NAND2_X1 U11118 ( .A1(s_IFID_IR[16]), .A2(s_IFID_IR[20]), .ZN(n19246) );
  NOR2_X1 U12081 ( .A1(n24616), .A2(n18059), .ZN(n20107) );
  NAND2_X1 U12043 ( .A1(s_IFID_IR[21]), .A2(n24610), .ZN(n20069) );
  NOR2_X1 U12038 ( .A1(s_IFID_IR[21]), .A2(n24610), .ZN(n20076) );
  NOR2_X1 U12016 ( .A1(n20069), .A2(n20080), .ZN(n19393) );
  NOR3_X1 U12201 ( .A1(s_IFID_IR[28]), .A2(n14191), .A3(n24583), .ZN(n19282)
         );
  AOI211_X1 U10648 ( .C1(n18312), .C2(n385), .A(n18740), .B(n18741), .ZN(
        n18733) );
  AOI22_X1 U10647 ( .A1(net716461), .A2(n377), .B1(n18347), .B2(n383), .ZN(
        n18734) );
  AOI22_X1 U10658 ( .A1(net767167), .A2(n374), .B1(n18326), .B2(n24758), .ZN(
        n18752) );
  AOI22_X1 U10657 ( .A1(n18300), .A2(n375), .B1(net767235), .B2(n24759), .ZN(
        n18744) );
  AOI22_X1 U10659 ( .A1(n18328), .A2(n17683), .B1(n18329), .B2(n17685), .ZN(
        n18751) );
  OAI22_X1 U10652 ( .A1(n399), .A2(n18315), .B1(n398), .B2(n18316), .ZN(n18740) );
  OAI211_X1 U10649 ( .C1(n391), .C2(net518461), .A(n18742), .B(n18743), .ZN(
        n18741) );
  AOI22_X1 U10654 ( .A1(n18307), .A2(n17687), .B1(net716405), .B2(n17686), 
        .ZN(n18747) );
  AOI22_X1 U10655 ( .A1(net767239), .A2(n24720), .B1(n18306), .B2(n386), .ZN(
        n18746) );
  AOI22_X1 U10656 ( .A1(n18310), .A2(n387), .B1(n18311), .B2(n373), .ZN(n18745) );
  AOI211_X1 U10643 ( .C1(n372), .C2(n18343), .A(n18737), .B(n18738), .ZN(
        n18736) );
  AOI22_X1 U10646 ( .A1(n18338), .A2(n381), .B1(n18339), .B2(n378), .ZN(n18735) );
  AOI22_X1 U10660 ( .A1(n18330), .A2(n379), .B1(n18331), .B2(n17684), .ZN(
        n18750) );
  AOI22_X1 U10651 ( .A1(net767173), .A2(n382), .B1(n18321), .B2(n384), .ZN(
        n18742) );
  NAND2_X1 U10650 ( .A1(n18529), .A2(n376), .ZN(n18743) );
  NOR2_X1 U10645 ( .A1(n397), .A2(net767232), .ZN(n18737) );
  OAI22_X1 U10644 ( .A1(n396), .A2(net767237), .B1(net716477), .B2(n24646), 
        .ZN(n18738) );
  AOI211_X1 U10803 ( .C1(n18312), .C2(n888), .A(n18933), .B(n18934), .ZN(
        n18926) );
  AOI22_X1 U10802 ( .A1(net716461), .A2(n880), .B1(n18347), .B2(n886), .ZN(
        n18927) );
  AOI22_X1 U10813 ( .A1(net767167), .A2(n877), .B1(n18326), .B2(n24752), .ZN(
        n18945) );
  AOI22_X1 U10812 ( .A1(n18300), .A2(n878), .B1(net767235), .B2(n24753), .ZN(
        n18937) );
  AOI22_X1 U10814 ( .A1(n18328), .A2(n17772), .B1(n18329), .B2(n17774), .ZN(
        n18944) );
  OAI22_X1 U10807 ( .A1(n902), .A2(n18315), .B1(n901), .B2(n18316), .ZN(n18933) );
  OAI211_X1 U10804 ( .C1(n894), .C2(net518461), .A(n18935), .B(n18936), .ZN(
        n18934) );
  AOI22_X1 U10809 ( .A1(n18307), .A2(n17776), .B1(net716405), .B2(n17775), 
        .ZN(n18940) );
  AOI22_X1 U10810 ( .A1(net767239), .A2(n24717), .B1(n18306), .B2(n889), .ZN(
        n18939) );
  AOI22_X1 U10811 ( .A1(n18310), .A2(n890), .B1(n18311), .B2(n876), .ZN(n18938) );
  AOI211_X1 U10798 ( .C1(n875), .C2(n18343), .A(n18930), .B(n18931), .ZN(
        n18929) );
  AOI22_X1 U10801 ( .A1(n18338), .A2(n884), .B1(n18339), .B2(n881), .ZN(n18928) );
  AOI22_X1 U10815 ( .A1(n18330), .A2(n882), .B1(n18331), .B2(n17773), .ZN(
        n18943) );
  AOI22_X1 U10806 ( .A1(net767173), .A2(n885), .B1(n18321), .B2(n887), .ZN(
        n18935) );
  NAND2_X1 U10805 ( .A1(n18529), .A2(n879), .ZN(n18936) );
  NOR2_X1 U10800 ( .A1(n900), .A2(net767232), .ZN(n18930) );
  OAI22_X1 U10799 ( .A1(n899), .A2(net767237), .B1(net716477), .B2(n24643), 
        .ZN(n18931) );
  SDFFR_X1 \core_inst/IDEX_IR/DFF_28/data_reg  ( .D(s_IFID_IR[28]), .SI(1'b0), 
        .SE(net796156), .CK(DLX_CLK), .RN(DLX_RST), .Q(n14073), .QN(net741237)
         );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_22/data_reg  ( .D(net712808), .SI(n23298), .SE(n22936), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [22]), .QN(net749434) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_15/data_reg  ( .D(n26530), 
        .SI(n24209), .SE(n22936), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [15]), .QN(n6516) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_27/data_reg  ( .D(n26559), 
        .SI(n24210), .SE(n24260), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [27]), .QN(n5171) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_17/data_reg  ( .D(n26534), 
        .SI(n24211), .SE(n24260), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [17]), .QN(n6511) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_30/data_reg  ( .D(n26410), 
        .SI(n24212), .SE(n22936), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/RES_GENERATOR/CSA_15/RCA_1/cout_tmp[0] ), .QN(n6546) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_5/data_reg  ( .D(n24263), 
        .SI(net734607), .SE(n24260), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [5]), .QN(n6514) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_25/data_reg  ( .D(n26458), 
        .SI(net749292), .SE(n22936), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [25]), .QN(n6402) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_24/data_reg  ( .D(n26571), 
        .SI(net754762), .SE(n24260), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [24]) );
  DFFRS_X1 \core_inst/IDEX_IMM_IN/DFF_18/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_18/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .QN(n23269) );
  DFFRS_X1 \core_inst/IDEX_IMM_IN/DFF_23/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_23/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .QN(n23264) );
  DFFRS_X1 \core_inst/IDEX_IMM_IN/DFF_21/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_21/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .QN(n23265) );
  DFFRS_X1 \core_inst/IDEX_IMM_IN/DFF_19/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_19/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .QN(n23267) );
  DFFRS_X1 \core_inst/IDEX_IMM_IN/DFF_20/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_20/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .QN(n23263) );
  DFFRS_X1 \core_inst/IDEX_IMM_IN/DFF_17/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_17/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .QN(n23268) );
  DFFRS_X1 \core_inst/IDEX_RF_IN2/DFF_21/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_21/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .QN(net780186) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_7/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_7/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        n25359) );
  DFFR_X1 \core_inst/IDEX_RF_IN1/DFF_12/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_12/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .QN(
        net740634) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_6/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_6/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n17667), .QN(n22699) );
  DFFRS_X1 \core_inst/IDEX_RF_IN2/DFF_3/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .QN(net780188) );
  DFFRS_X1 \core_inst/IDEX_RF_IN1/DFF_6/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_6/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .Q(n25342) );
  DFFRS_X1 \core_inst/IDEX_RF_IN1/DFF_5/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_5/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .Q(net399701) );
  DFFRS_X1 \core_inst/IDEX_RF_IN1/DFF_2/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_2/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .Q(n17664) );
  DFFRS_X1 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_1/data_reg  ( .D(
        \core_inst/IF_stage/PROGRAM_COUNTER/DFF_1/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .SN(1'b1), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [1]) );
  AOI22_X1 U11785 ( .A1(n19336), .A2(n24712), .B1(n19337), .B2(n17814), .ZN(
        n19905) );
  AOI22_X1 U11788 ( .A1(n19372), .A2(n17820), .B1(n19373), .B2(n17819), .ZN(
        n19910) );
  NOR4_X1 U11775 ( .A1(n19901), .A2(n19902), .A3(n19903), .A4(n19904), .ZN(
        n19895) );
  AOI22_X1 U11773 ( .A1(n19308), .A2(n24714), .B1(n23995), .B2(n17822), .ZN(
        n19896) );
  OAI22_X1 U11779 ( .A1(n2883), .A2(n19350), .B1(n2882), .B2(n26614), .ZN(
        n19901) );
  OAI22_X1 U11778 ( .A1(n2873), .A2(n19396), .B1(n25677), .B2(n24639), .ZN(
        n19902) );
  OAI22_X1 U11777 ( .A1(n2880), .A2(n25678), .B1(n25676), .B2(n24640), .ZN(
        n19903) );
  OAI22_X1 U11776 ( .A1(n2879), .A2(n19370), .B1(n2877), .B2(n19365), .ZN(
        n19904) );
  AOI22_X1 U11781 ( .A1(n24026), .A2(n24713), .B1(n19333), .B2(n17811), .ZN(
        n19908) );
  AOI22_X1 U11783 ( .A1(n25674), .A2(n17809), .B1(n25680), .B2(n17815), .ZN(
        n19907) );
  AOI22_X1 U11784 ( .A1(n24007), .A2(n17813), .B1(n19335), .B2(n17816), .ZN(
        n19906) );
  AOI211_X1 U11769 ( .C1(n23994), .C2(n17810), .A(n19899), .B(n19900), .ZN(
        n19898) );
  AOI22_X1 U11772 ( .A1(n19315), .A2(n17823), .B1(n25683), .B2(n17821), .ZN(
        n19897) );
  NOR2_X1 U11771 ( .A1(n2892), .A2(n19389), .ZN(n19899) );
  OAI22_X1 U11770 ( .A1(n2896), .A2(n19378), .B1(n2895), .B2(n19388), .ZN(
        n19900) );
  DFFRS_X1 \core_inst/IDEX_RF_IN1/DFF_15/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_15/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .QN(n23266) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_18/data_reg  ( .D(net713438), .SI(n24099), .SE(net826165), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [18]) );
  AOI22_X1 U11892 ( .A1(n19336), .A2(n24704), .B1(n19337), .B2(n17865), .ZN(
        n19989) );
  AOI22_X1 U11895 ( .A1(n19372), .A2(n17871), .B1(n19373), .B2(n17870), .ZN(
        n19994) );
  NOR4_X1 U11882 ( .A1(n19985), .A2(n19986), .A3(n19987), .A4(n19988), .ZN(
        n19979) );
  AOI22_X1 U11880 ( .A1(n19308), .A2(n24706), .B1(n23995), .B2(n17873), .ZN(
        n19980) );
  OAI22_X1 U11886 ( .A1(n3027), .A2(n19350), .B1(n3026), .B2(n26614), .ZN(
        n19985) );
  OAI22_X1 U11885 ( .A1(n3017), .A2(n19396), .B1(n25677), .B2(n24633), .ZN(
        n19986) );
  OAI22_X1 U11884 ( .A1(n3024), .A2(n25678), .B1(n25676), .B2(n24634), .ZN(
        n19987) );
  OAI22_X1 U11883 ( .A1(n3023), .A2(n19370), .B1(n3021), .B2(n19365), .ZN(
        n19988) );
  AOI22_X1 U11888 ( .A1(n19332), .A2(n24705), .B1(n25682), .B2(n17862), .ZN(
        n19992) );
  AOI22_X1 U11890 ( .A1(n25674), .A2(n17860), .B1(n25680), .B2(n17866), .ZN(
        n19991) );
  AOI22_X1 U11891 ( .A1(n24007), .A2(n17864), .B1(n19335), .B2(n17867), .ZN(
        n19990) );
  AOI211_X1 U11876 ( .C1(n23994), .C2(n17861), .A(n19983), .B(n19984), .ZN(
        n19982) );
  AOI22_X1 U11879 ( .A1(n19315), .A2(n17874), .B1(n25683), .B2(n17872), .ZN(
        n19981) );
  NOR2_X1 U11878 ( .A1(n3036), .A2(n19389), .ZN(n19983) );
  OAI22_X1 U11877 ( .A1(n3040), .A2(n19378), .B1(n3039), .B2(n19388), .ZN(
        n19984) );
  AOI22_X1 U11944 ( .A1(n19336), .A2(n24698), .B1(n19337), .B2(n18009), .ZN(
        n20031) );
  AOI22_X1 U11947 ( .A1(n19372), .A2(n18015), .B1(n19373), .B2(n18014), .ZN(
        n20036) );
  NOR4_X1 U11934 ( .A1(n20027), .A2(n20028), .A3(n20029), .A4(n20030), .ZN(
        n20021) );
  AOI22_X1 U11932 ( .A1(n19308), .A2(n24700), .B1(n23995), .B2(n18017), .ZN(
        n20022) );
  OAI22_X1 U11938 ( .A1(n2703), .A2(n19350), .B1(n2702), .B2(n26614), .ZN(
        n20027) );
  OAI22_X1 U11937 ( .A1(n2693), .A2(n19396), .B1(n25677), .B2(n24629), .ZN(
        n20028) );
  OAI22_X1 U11936 ( .A1(n2700), .A2(n25678), .B1(n25676), .B2(n24630), .ZN(
        n20029) );
  OAI22_X1 U11935 ( .A1(n2699), .A2(n19370), .B1(n2697), .B2(n19365), .ZN(
        n20030) );
  AOI22_X1 U11940 ( .A1(n19332), .A2(n24699), .B1(n25682), .B2(n18006), .ZN(
        n20034) );
  AOI22_X1 U11942 ( .A1(n25674), .A2(n18004), .B1(n25680), .B2(n18010), .ZN(
        n20033) );
  AOI22_X1 U11943 ( .A1(n24007), .A2(n18008), .B1(n19335), .B2(n18011), .ZN(
        n20032) );
  AOI211_X1 U11928 ( .C1(n23994), .C2(n18005), .A(n20025), .B(n20026), .ZN(
        n20024) );
  AOI22_X1 U11931 ( .A1(n19315), .A2(n18018), .B1(n25683), .B2(n18016), .ZN(
        n20023) );
  NOR2_X1 U11930 ( .A1(n2712), .A2(n19389), .ZN(n20025) );
  OAI22_X1 U11929 ( .A1(n2716), .A2(n19378), .B1(n2715), .B2(n19388), .ZN(
        n20026) );
  DFFRS_X1 \core_inst/IDEX_RF_IN1/DFF_1/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .Q(n14764) );
  NOR2_X1 U11121 ( .A1(s_IFID_IR[16]), .A2(net741525), .ZN(n19255) );
  NOR2_X1 U12084 ( .A1(n14210), .A2(n24677), .ZN(n20110) );
  NOR2_X1 U12019 ( .A1(n20081), .A2(n20068), .ZN(n19334) );
  INV_X1 U12008 ( .A(n20071), .ZN(n20067) );
  INV_X1 U11094 ( .A(n19250), .ZN(n19245) );
  NAND3_X1 U15903 ( .A1(n19288), .A2(s_ID_rf_write_en), .A3(n19291), .ZN(
        n20200) );
  INV_X1 U12003 ( .A(n20061), .ZN(n20066) );
  INV_X1 U12080 ( .A(n20107), .ZN(n20111) );
  INV_X1 U11995 ( .A(n20080), .ZN(n20060) );
  INV_X1 U12042 ( .A(n20069), .ZN(n20062) );
  INV_X1 U12082 ( .A(n20110), .ZN(n18188) );
  INV_X1 U12015 ( .A(n20070), .ZN(n20064) );
  INV_X1 U12034 ( .A(n20068), .ZN(n20078) );
  INV_X1 U11089 ( .A(n19239), .ZN(n19244) );
  INV_X1 U11090 ( .A(n19265), .ZN(n19264) );
  INV_X1 U11081 ( .A(n19261), .ZN(n19238) );
  INV_X1 U11125 ( .A(n19248), .ZN(n19240) );
  INV_X1 U13810 ( .A(n19288), .ZN(n20396) );
  INV_X1 U13503 ( .A(n19291), .ZN(n20397) );
  INV_X1 U11117 ( .A(n19246), .ZN(n19257) );
  INV_X1 U11100 ( .A(n19249), .ZN(n19242) );
  NAND3_X1 U15904 ( .A1(n19289), .A2(n19292), .A3(n26780), .ZN(n20153) );
  NAND3_X1 U15897 ( .A1(n19294), .A2(n20609), .A3(n20610), .ZN(n20220) );
  NAND3_X1 U15901 ( .A1(n19294), .A2(n19289), .A3(n20610), .ZN(n20372) );
  INV_X1 U11082 ( .A(n18343), .ZN(n18401) );
  NAND3_X1 U15898 ( .A1(n19292), .A2(n20609), .A3(n26780), .ZN(n20240) );
  NAND3_X1 U15900 ( .A1(n19289), .A2(n26780), .A3(n20610), .ZN(n20332) );
  NAND3_X1 U15899 ( .A1(n19294), .A2(n19292), .A3(n20609), .ZN(n20260) );
  INV_X1 U11751 ( .A(n19372), .ZN(n19323) );
  NAND4_X1 U10201 ( .A1(s_MEM_LOAD_TYPE[1]), .A2(s_MEM_SIGNED_LOAD), .A3(
        \core_inst/MEM/MUX_LOAD/MUX_BIT_7/s_top ), .A4(n24774), .ZN(n18198) );
  INV_X1 U11996 ( .A(n19348), .ZN(n19396) );
  NAND3_X1 U15896 ( .A1(n20609), .A2(n26780), .A3(n20610), .ZN(n20201) );
  INV_X1 U11739 ( .A(n19365), .ZN(n19345) );
  INV_X1 U11747 ( .A(n19395), .ZN(n19327) );
  INV_X1 U11750 ( .A(n19373), .ZN(n19324) );
  INV_X1 U11740 ( .A(n19370), .ZN(n19344) );
  INV_X1 U11825 ( .A(n19389), .ZN(n19314) );
  INV_X1 U11752 ( .A(n19383), .ZN(n19320) );
  INV_X1 U10133 ( .A(n26777), .ZN(n18139) );
  INV_X1 U12032 ( .A(n19326), .ZN(n19530) );
  INV_X1 U11829 ( .A(n19378), .ZN(n19318) );
  INV_X1 U11827 ( .A(n19388), .ZN(n19319) );
  INV_X1 U10141 ( .A(n18193), .ZN(n18151) );
  NOR2_X1 U13941 ( .A1(n18046), .A2(n18039), .ZN(n19292) );
  NOR2_X1 U13940 ( .A1(n18046), .A2(n18038), .ZN(n19294) );
  NOR2_X1 U13942 ( .A1(n18046), .A2(n18040), .ZN(n19289) );
  NOR2_X1 U13937 ( .A1(n18046), .A2(n18042), .ZN(n19291) );
  NOR2_X1 U13938 ( .A1(n18046), .A2(n18041), .ZN(n19288) );
  INV_X1 U13707 ( .A(n19289), .ZN(n20609) );
  INV_X1 U13809 ( .A(n19292), .ZN(n20610) );
  NAND3_X1 U15902 ( .A1(s_ID_rf_write_en), .A2(n19291), .A3(n20396), .ZN(
        n20154) );
  NAND3_X1 U15893 ( .A1(s_ID_rf_write_en), .A2(n20396), .A3(n20397), .ZN(
        n20293) );
  NAND3_X1 U15894 ( .A1(s_ID_rf_write_en), .A2(n19288), .A3(n20397), .ZN(
        n20431) );
  INV_X1 U11978 ( .A(n19384), .ZN(n19315) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_4/data_reg  ( .D(n26605), 
        .SI(n24128), .SE(net812941), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [4]) );
  DFFR_X1 \cu_inst/EX/DFF_16/data_reg  ( .D(\cu_inst/EX/DFF_16/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(net366531), .QN(net741456) );
  DFFR_X1 \core_inst/IFID_IR/DFF_3/data_reg  ( .D(\core_inst/IFID_IR/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n14128), .QN(n24585) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_24/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_24/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_24/N3 ), .QN(n6740) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_19/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_19/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_19/N3 ), .QN(n13805) );
  DFFR_X1 \core_inst/IFID_IR/DFF_1/data_reg  ( .D(\core_inst/IFID_IR/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n18059) );
  DFFR_X1 \core_inst/IFID_IR/DFF_30/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_30/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_IFID_IR[30]), .QN(net741565) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_11/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_11/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_11/N3 ), .QN(n1182) );
  DFFR_X1 \core_inst/IFID_IR/DFF_29/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_29/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_IFID_IR[29]), .QN(n24583) );
  DFFR_X1 \core_inst/IFID_IR/DFF_27/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_27/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_IFID_IR[27]), .QN(n24581) );
  DFFR_X1 \core_inst/IFID_IR/DFF_13/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_13/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n25336)
         );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_31/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_31/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_31/N3 ), .QN(n478) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_17/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_17/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_17/N3 ), .QN(n17743) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_5/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_5/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_5/N3 ), .QN(n1378) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_22/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_22/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_22/N3 ), .QN(n829) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_20/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_20/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_20/N3 ), .QN(n869) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_16/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_16/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_16/N3 ), .QN(n5585) );
  DFFR_X1 \core_inst/EXMEM_IR/DFF_11/data_reg  ( .D(
        \core_inst/EXMEM_IR/DFF_11/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_IR/DFF_11/N3 ), .QN(n5181) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_20/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_20/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_20/N3 ), .QN(n1702) );
  DFFR_X1 \core_inst/IFID_IR/DFF_0/data_reg  ( .D(\core_inst/IFID_IR/DFF_0/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n14190), .QN(n24680) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_4/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_4/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_4/N3 ), .QN(n1704) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_8/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_8/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_8/N3 ), .QN(n1726) );
  DFFR_X1 \core_inst/IFID_IR/DFF_22/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_22/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_IFID_IR[22]), .QN(n24618) );
  DFFR_X1 \core_inst/IFID_IR/DFF_28/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_28/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_IFID_IR[28]), .QN(n24611) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_3/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_3/N3 ), .QN(n1456) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_12/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_12/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_12/N3 ), .QN(n1744) );
  DFFR_X1 \core_inst/IFID_IR/DFF_16/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_16/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_IFID_IR[16]), .QN(n24527) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_15/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_15/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_15/N3 ), .QN(n1064) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_8/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_8/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_8/N3 ), .QN(n5582) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_28/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_28/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_28/N3 ), .QN(n1716) );
  DFFR_X1 \core_inst/IFID_IR/DFF_26/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_26/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_IFID_IR[26]), .QN(n24584) );
  DFFR_X1 \core_inst/IFID_IR/DFF_25/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_25/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_IFID_IR[25]), .QN(n24610) );
  DFFR_X1 \core_inst/EXMEM_IR/DFF_26/data_reg  ( .D(
        \core_inst/EXMEM_IR/DFF_26/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(n14429), .QN(n17659) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_21/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_21/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_21/N3 ), .QN(n1698) );
  DFFR_X1 \core_inst/EXMEM_IR/DFF_12/data_reg  ( .D(
        \core_inst/EXMEM_IR/DFF_12/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_IR/DFF_12/N3 ), .QN(n1637) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_1/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        net741280), .QN(n1501) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_0/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_0/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n25334), .QN(n1539) );
  DFFR_X1 \core_inst/EXMEM_IR/DFF_17/data_reg  ( .D(
        \core_inst/EXMEM_IR/DFF_17/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_IR/DFF_17/N3 ), .QN(n5174) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_22/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_22/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_22/N3 ), .QN(n1736) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_17/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_17/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_17/N3 ), .QN(n1740) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_24/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_24/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_24/N3 ), .QN(n1720) );
  DFFR_X1 \core_inst/EXMEM_IR/DFF_16/data_reg  ( .D(
        \core_inst/EXMEM_IR/DFF_16/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_IR/DFF_16/N3 ), .QN(n5598) );
  DFFR_X1 \core_inst/EXMEM_IR/DFF_13/data_reg  ( .D(
        \core_inst/EXMEM_IR/DFF_13/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_IR/DFF_13/N3 ), .QN(n5607) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_31/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_31/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_31/N3 ), .QN(n1752) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_21/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_21/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_21/N3 ), .QN(n5587) );
  DFFR_X1 \core_inst/EXMEM_IR/DFF_20/data_reg  ( .D(
        \core_inst/EXMEM_IR/DFF_20/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_IR/DFF_20/N3 ), .QN(n5613) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_5/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_5/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_5/N3 ), .QN(n1694) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_25/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_25/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_25/N3 ), .QN(net81266) );
  DFFR_X1 \core_inst/IDEX_NPC/DFF_9/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_9/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_9/N3 ), .QN(n367) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_27/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_27/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_27/N3 ), .QN(n1742) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_25/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_25/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_25/N3 ), .QN(n1738) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_3/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_3/N3 ), .QN(n1692) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_19/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_19/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_19/N3 ), .QN(n1718) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_16/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_16/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_16/N3 ), .QN(n1708) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_10/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_10/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_10/N3 ), .QN(n1748) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_18/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_18/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_18/N3 ), .QN(n1722) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_9/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_9/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_9/N3 ), .QN(n1714) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_11/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_11/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_11/N3 ), .QN(n1746) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_7/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_7/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_7/N3 ), .QN(n1696) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_15/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_15/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_15/N3 ), .QN(n1710) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_29/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_29/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_29/N3 ), .QN(n1730) );
  DFFR_X1 \core_inst/EXMEM_ALU_OUT/DFF_0/data_reg  ( .D(
        \core_inst/EXMEM_ALU_OUT/DFF_0/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/MEMWB_ALUOUT/DFF_0/N3 ), .QN(n1750) );
  DFFS_X1 \core_inst/EXMEM_DATAIN/DFF_9/data_reg  ( .D(n23946), .CK(DLX_CLK), 
        .SN(DLX_RST), .QN(\core_inst/ps_EXMEM_DATA_IN [9]) );
  SDFFR_X2 \core_inst/IFID_IR/DFF_2/data_reg  ( .D(
        \core_inst/s_IF_OUT_IR_OUT [2]), .SI(1'b0), .SE(net796200), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(n14195), .QN(n24616) );
  DFFS_X1 \core_inst/EXMEM_IR/DFF_31/data_reg  ( .D(
        \core_inst/EXMEM_IR/DFF_31/data_reg/n15 ), .CK(DLX_CLK), .SN(DLX_RST), 
        .Q(net741339), .QN(net89524) );
  NAND2_X1 U10160 ( .A1(n18201), .A2(n18206), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_28/N3 ) );
  NAND2_X1 U10179 ( .A1(n18201), .A2(n18215), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_19/N3 ) );
  NAND2_X1 U10172 ( .A1(n18201), .A2(n18212), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_22/N3 ) );
  NAND2_X1 U10183 ( .A1(n18201), .A2(n18217), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_17/N3 ) );
  NAND2_X1 U10168 ( .A1(n18201), .A2(n18210), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_24/N3 ) );
  NAND2_X1 U10176 ( .A1(n18201), .A2(n18214), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_20/N3 ) );
  NAND2_X1 U10155 ( .A1(n18201), .A2(n18204), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_30/N3 ) );
  NAND2_X1 U10164 ( .A1(n18201), .A2(n18208), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_26/N3 ) );
  NAND2_X1 U10153 ( .A1(n18201), .A2(n18202), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_31/N3 ) );
  NAND2_X1 U10185 ( .A1(n18201), .A2(n18218), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_16/N3 ) );
  OAI21_X1 U10190 ( .B1(s_MEM_LOAD_TYPE[1]), .B2(n18220), .A(n18198), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_15/N3 ) );
  NAND2_X1 U10166 ( .A1(n18201), .A2(n18209), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_25/N3 ) );
  NAND2_X1 U10174 ( .A1(n18201), .A2(n18213), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_21/N3 ) );
  NAND2_X1 U10162 ( .A1(n18201), .A2(n18207), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_27/N3 ) );
  NAND2_X1 U10170 ( .A1(n18201), .A2(n18211), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_23/N3 ) );
  NAND2_X1 U10181 ( .A1(n18201), .A2(n18216), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_18/N3 ) );
  NAND2_X1 U10158 ( .A1(n18201), .A2(n18205), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_29/N3 ) );
  NOR2_X1 U12074 ( .A1(n18062), .A2(n14128), .ZN(n20108) );
  AOI21_X1 U12070 ( .B1(n20108), .B2(n18161), .A(n18146), .ZN(n18169) );
  NAND2_X1 U12083 ( .A1(n20110), .A2(n24585), .ZN(n20113) );
  OAI21_X1 U12076 ( .B1(n14195), .B2(n20113), .A(n18140), .ZN(n18150) );
  NOR3_X1 U12193 ( .A1(s_IFID_IR[27]), .A2(n24611), .A3(n24583), .ZN(n20133)
         );
  OAI21_X1 U10200 ( .B1(s_MEM_LOAD_TYPE[1]), .B2(n18225), .A(n18198), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_10/N3 ) );
  OAI21_X1 U10147 ( .B1(s_MEM_LOAD_TYPE[1]), .B2(n18199), .A(n18198), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_8/N3 ) );
  OAI21_X1 U10145 ( .B1(s_MEM_LOAD_TYPE[1]), .B2(n18197), .A(n18198), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_9/N3 ) );
  OAI21_X1 U10198 ( .B1(s_MEM_LOAD_TYPE[1]), .B2(n18224), .A(n18198), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_11/N3 ) );
  OAI21_X1 U10192 ( .B1(s_MEM_LOAD_TYPE[1]), .B2(n18221), .A(n18198), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_14/N3 ) );
  OAI21_X1 U10194 ( .B1(s_MEM_LOAD_TYPE[1]), .B2(n18222), .A(n18198), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_13/N3 ) );
  OAI21_X1 U10196 ( .B1(s_MEM_LOAD_TYPE[1]), .B2(n18223), .A(n18198), .ZN(
        \core_inst/MEMWB_DATAOUT/DFF_12/N3 ) );
  NAND3_X1 U15843 ( .A1(n18171), .A2(n26779), .A3(n18172), .ZN(n18167) );
  AOI221_X1 U10124 ( .B1(n14190), .B2(n18169), .C1(n18170), .C2(n18169), .A(
        n18139), .ZN(n18168) );
  AOI21_X1 U10123 ( .B1(n18166), .B2(n18167), .A(n18168), .ZN(n18165) );
  NAND2_X1 U10122 ( .A1(n18164), .A2(n18165), .ZN(\cu_inst/EX/DFF_14/N3 ) );
  OAI211_X1 U10121 ( .C1(n18161), .C2(n18162), .A(n26777), .B(n24585), .ZN(
        n18160) );
  OAI221_X1 U10120 ( .B1(n24584), .B2(n18158), .C1(n24584), .C2(n18159), .A(
        n18160), .ZN(n18157) );
  AOI21_X1 U10119 ( .B1(n18145), .B2(n18156), .A(n18157), .ZN(n18155) );
  OAI211_X1 U10118 ( .C1(s_IFID_IR[30]), .C2(n18153), .A(n18154), .B(n18155), 
        .ZN(\cu_inst/EX/DFF_15/N3 ) );
  DFFR_X2 \cu_inst/EX/DFF_11/data_reg  ( .D(\cu_inst/EX/DFF_11/N3 ), .CK(
        DLX_CLK), .RN(DLX_RST), .Q(net741726), .QN(net741686) );
  DFFR_X1 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_12/data_reg  ( .D(n26782), 
        .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [12]), .QN(n24343) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_19/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_19/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n22941), .QN(n874) );
  DFFRS_X1 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_16/data_reg  ( .D(n16384), 
        .CK(DLX_CLK), .RN(DLX_RST), .SN(1'b1), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [16]) );
  DFFS_X1 \core_inst/IDEX_RF_IN1/DFF_16/data_reg  ( .D(n26328), .CK(DLX_CLK), 
        .SN(DLX_RST), .Q(n25361) );
  DFFS_X1 \core_inst/IDEX_RF_IN1/DFF_31/data_reg  ( .D(n26362), .CK(DLX_CLK), 
        .SN(DLX_RST), .Q(n25362) );
  DFFS_X1 \core_inst/IDEX_RF_IN2/DFF_9/data_reg  ( .D(n26685), .CK(DLX_CLK), 
        .SN(DLX_RST), .Q(n5610), .QN(n22816) );
  DFFS_X1 \core_inst/IDEX_RF_IN1/DFF_18/data_reg  ( .D(n26638), .CK(DLX_CLK), 
        .SN(DLX_RST), .Q(n25356) );
  DFFS_X1 \core_inst/IDEX_RF_IN2/DFF_15/data_reg  ( .D(n26651), .CK(DLX_CLK), 
        .SN(DLX_RST), .Q(n25324), .QN(n22944) );
  DFFS_X1 \core_inst/IDEX_RF_IN2/DFF_12/data_reg  ( .D(n26696), .CK(DLX_CLK), 
        .SN(DLX_RST), .Q(n5611) );
  DFFS_X1 \core_inst/IDEX_RF_IN2/DFF_11/data_reg  ( .D(n26302), .CK(DLX_CLK), 
        .SN(DLX_RST), .Q(n25325), .QN(n22943) );
  DFFS_X1 \core_inst/IDEX_RF_IN1/DFF_17/data_reg  ( .D(n26403), .CK(DLX_CLK), 
        .SN(DLX_RST), .Q(n25364) );
  DFFS_X1 \core_inst/IDEX_IMM_IN/DFF_25/data_reg  ( .D(n23944), .CK(DLX_CLK), 
        .SN(DLX_RST), .QN(n14464) );
  DFFS_X1 \core_inst/IDEX_RF_IN1/DFF_26/data_reg  ( .D(n26333), .CK(DLX_CLK), 
        .SN(DLX_RST), .QN(n25341) );
  DFFS_X1 \core_inst/IDEX_RF_IN1/DFF_28/data_reg  ( .D(n26392), .CK(DLX_CLK), 
        .SN(DLX_RST), .QN(n14758) );
  DFFS_X1 \core_inst/IDEX_RF_IN1/DFF_30/data_reg  ( .D(n26312), .CK(DLX_CLK), 
        .SN(DLX_RST), .QN(n25343) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_28/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_28/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n25332), .QN(n5602) );
  DFFR_X1 \core_inst/IFID_IR/DFF_20/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_20/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_IFID_IR[20]), .QN(net741525) );
  DFFS_X1 \core_inst/IDEX_RF_IN1/DFF_25/data_reg  ( .D(n26470), .CK(DLX_CLK), 
        .SN(DLX_RST), .QN(n25353) );
  DFFRS_X1 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_0/data_reg  ( .D(
        \core_inst/IF_stage/PROGRAM_COUNTER/DFF_0/N3 ), .CK(DLX_CLK), .RN(
        DLX_RST), .SN(1'b1), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/CLA_PG_NET/N1 ) );
  DFFRS_X1 \core_inst/IDEX_RF_IN2/DFF_30/data_reg  ( .D(n22714), .CK(DLX_CLK), 
        .RN(DLX_RST), .SN(1'b1), .Q(n22855), .QN(n22672) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_20/data_reg  ( .D(net712793), .SI(n22856), .SE(net716331), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [20]), .QN(net749439) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_21/data_reg  ( .D(n22866), 
        .SI(net794712), .SE(net796271), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [21]), .QN(n6461) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_25/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_25/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n25331), .QN(n371) );
  DFFR_X1 \core_inst/IDEX_RF_IN2/DFF_17/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_17/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        n22814), .QN(n680) );
  DFFRS_X1 \core_inst/IDEX_RF_IN2/DFF_18/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_18/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .QN(n22676) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_23/data_reg  ( .D(n26257), 
        .SI(n24123), .SE(net796271), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [23]), .QN(n6462) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_31/data_reg  ( .D(n25446), 
        .SI(n22682), .SE(net716331), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/RES_GENERATOR/CSA_15/sum_rca_0[1] ) );
  DFFRS_X1 \core_inst/IDEX_RF_IN2/DFF_26/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_26/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .QN(n22677) );
  DFFR_X1 \core_inst/IFID_IR/DFF_23/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_23/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_IFID_IR[23]), .QN(n24582) );
  DFFRS_X1 \core_inst/IDEX_IMM_IN/DFF_24/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_24/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .QN(n23271) );
  NAND2_X1 U10108 ( .A1(n18130), .A2(n18131), .ZN(\cu_inst/EX/DFF_7/N3 ) );
  NOR3_X1 U10140 ( .A1(net741279), .A2(n18151), .A3(n18137), .ZN(n18131) );
  OR2_X1 U10112 ( .A1(n18136), .A2(n18137), .ZN(\cu_inst/EX/DFF_3/N3 ) );
  NAND3_X1 U15866 ( .A1(net741620), .A2(net741547), .A3(net741696), .ZN(n19262) );
  NAND3_X1 U15865 ( .A1(s_IFID_IR[18]), .A2(s_IFID_IR[19]), .A3(net741620), 
        .ZN(n19243) );
  NOR3_X1 U11127 ( .A1(s_IFID_IR[18]), .A2(s_IFID_IR[19]), .A3(net741620), 
        .ZN(n19265) );
  NOR3_X1 U11095 ( .A1(net741620), .A2(net741547), .A3(net741696), .ZN(n19250)
         );
  DFFRS_X1 \core_inst/IDEX_IMM_IN/DFF_27/data_reg  ( .D(n24573), .CK(DLX_CLK), 
        .RN(DLX_RST), .SN(1'b1), .QN(n22687) );
  DFFRS_X1 \core_inst/IDEX_IMM_IN/DFF_31/data_reg  ( .D(n24573), .CK(DLX_CLK), 
        .RN(DLX_RST), .SN(1'b1), .Q(n25345) );
  DFFRS_X1 \core_inst/IDEX_IMM_IN/DFF_26/data_reg  ( .D(n24573), .CK(DLX_CLK), 
        .RN(DLX_RST), .SN(1'b1), .QN(n6156) );
  DFFRS_X1 \core_inst/IDEX_IMM_IN/DFF_30/data_reg  ( .D(n6695), .CK(DLX_CLK), 
        .RN(DLX_RST), .SN(1'b1), .QN(n22688) );
  DFFRS_X1 \core_inst/IDEX_IMM_IN/DFF_28/data_reg  ( .D(n6695), .CK(DLX_CLK), 
        .RN(DLX_RST), .SN(1'b1), .Q(n17674) );
  DFFRS_X1 \core_inst/IDEX_IMM_IN/DFF_29/data_reg  ( .D(n6695), .CK(DLX_CLK), 
        .RN(DLX_RST), .SN(1'b1), .Q(n17675) );
  DFFRS_X1 \core_inst/IDEX_RF_IN1/DFF_11/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_11/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .QN(n22686) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_14/data_reg  ( .D(net712486), .SI(n22759), .SE(net716331), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [14]) );
  DFFRS_X1 \core_inst/EXMEM_DATAIN/DFF_31/data_reg  ( .D(
        \core_inst/EXMEM_DATAIN/DFF_31/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .Q(\core_inst/ps_EXMEM_DATA_IN [31]) );
  DFFRS_X1 \core_inst/EXMEM_RF_ADDR_DEST/DFF_3/data_reg  ( .D(
        \core_inst/EXMEM_RF_ADDR_DEST/DFF_3/N3 ), .CK(DLX_CLK), .RN(DLX_RST), 
        .SN(1'b1), .Q(\core_inst/MEMWB_RF_ADDR_DEST/DFF_3/N3 ) );
  DFFRS_X1 \core_inst/IDEX_NPC/DFF_30/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_30/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(1'b1), 
        .Q(\core_inst/EXMEM_NPC/DFF_30/N3 ) );
  DFFRS_X1 \core_inst/IDEX_NPC/DFF_26/data_reg  ( .D(
        \core_inst/IDEX_NPC/DFF_26/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(1'b1), 
        .Q(\core_inst/EXMEM_NPC/DFF_26/N3 ) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_6/data_reg  ( .D(n24168), 
        .SI(n24134), .SE(net812284), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [6]) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_8/data_reg  ( .D(n23938), 
        .SI(n22745), .SE(net742593), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [8]) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_29/data_reg  ( .D(n26568), 
        .SI(n22940), .SE(net812284), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [29]), .QN(n6180) );
  SDFFR_X2 \core_inst/IDEX_NPC/DFF_23/data_reg  ( .D(n17757), .SI(1'b0), .SE(
        net826165), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/EXMEM_NPC/DFF_23/N3 ), .QN(n790) );
  DFFRS_X1 \core_inst/IDEX_IMM_IN/DFF_22/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_22/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .QN(n23270) );
  DFFRS_X1 \core_inst/IDEX_RF_ADDR_DEST/DFF_1/data_reg  ( .D(
        \core_inst/IDEX_RF_ADDR_DEST/DFF_1/N3 ), .CK(DLX_CLK), .RN(DLX_RST), 
        .SN(1'b1), .QN(n22811) );
  DFFRS_X1 \core_inst/IDEX_IMM_IN/DFF_16/data_reg  ( .D(
        \core_inst/IDEX_IMM_IN/DFF_16/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .Q(n25344) );
  DFFR_X1 \core_inst/IFID_IR/DFF_19/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_19/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_IFID_IR[19]), .QN(net741696) );
  AOI22_X1 U10725 ( .A1(n18328), .A2(n17758), .B1(n18329), .B2(n17760), .ZN(
        n18832) );
  AOI22_X1 U10723 ( .A1(n18300), .A2(n799), .B1(net767235), .B2(net741384), 
        .ZN(n18825) );
  AOI22_X1 U10724 ( .A1(net767167), .A2(n798), .B1(net716417), .B2(net741385), 
        .ZN(n18833) );
  AOI22_X1 U10726 ( .A1(n18330), .A2(n803), .B1(n18331), .B2(n17759), .ZN(
        n18831) );
  AOI22_X1 U10712 ( .A1(n18338), .A2(n805), .B1(n18339), .B2(n802), .ZN(n18816) );
  OAI22_X1 U10710 ( .A1(n820), .A2(net767237), .B1(net716477), .B2(net741518), 
        .ZN(n18819) );
  NOR2_X1 U10711 ( .A1(n821), .A2(net767232), .ZN(n18818) );
  AOI211_X1 U10709 ( .C1(n796), .C2(n18343), .A(n18818), .B(n18819), .ZN(
        n18817) );
  AOI22_X1 U10713 ( .A1(net716461), .A2(n801), .B1(n18347), .B2(n807), .ZN(
        n18815) );
  AOI22_X1 U10722 ( .A1(n18310), .A2(n811), .B1(n18311), .B2(n797), .ZN(n18826) );
  AOI22_X1 U10721 ( .A1(net767239), .A2(net741440), .B1(n18306), .B2(n810), 
        .ZN(n18827) );
  AOI22_X1 U10720 ( .A1(n18307), .A2(n17762), .B1(net716405), .B2(n17761), 
        .ZN(n18828) );
  NAND2_X1 U10716 ( .A1(n18529), .A2(n800), .ZN(n18824) );
  AOI22_X1 U10717 ( .A1(net767173), .A2(n806), .B1(n18321), .B2(n808), .ZN(
        n18823) );
  OAI211_X1 U10715 ( .C1(n815), .C2(net518461), .A(n18823), .B(n18824), .ZN(
        n18822) );
  OAI22_X1 U10718 ( .A1(n823), .A2(n18315), .B1(n822), .B2(n18316), .ZN(n18821) );
  AOI211_X1 U10714 ( .C1(n18312), .C2(n809), .A(n18821), .B(n18822), .ZN(
        n18814) );
  SDFFR_X2 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_3/data_reg  ( .D(n25580), 
        .SI(n26744), .SE(net716253), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_up_network_p[1] ), .QN(n6746) );
  DFFRS_X1 \core_inst/IDEX_RF_IN1/DFF_14/data_reg  ( .D(
        \core_inst/IDEX_RF_IN1/DFF_14/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .Q(n11928) );
  DFFR_X1 \core_inst/IFID_IR/DFF_18/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_18/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_IFID_IR[18]), .QN(net741547) );
  DFFR_X1 \core_inst/IFID_IR/DFF_24/data_reg  ( .D(
        \core_inst/IFID_IR/DFF_24/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .Q(
        s_IFID_IR[24]), .QN(n24586) );
  DFFRS_X1 \core_inst/IF_stage/PROGRAM_COUNTER/DFF_28/data_reg  ( .D(net521855), .CK(DLX_CLK), .RN(DLX_RST), .SN(1'b1), .Q(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [28]) );
  DFFRS_X1 \core_inst/IDEX_RF_IN2/DFF_20/data_reg  ( .D(
        \core_inst/IDEX_RF_IN2/DFF_20/N3 ), .CK(DLX_CLK), .RN(DLX_RST), .SN(
        1'b1), .Q(n22669) );
  NOR2_X1 U11103 ( .A1(n19249), .A2(n19246), .ZN(n18329) );
  AOI22_X1 U10769 ( .A1(n18328), .A2(n17765), .B1(n18329), .B2(n17767), .ZN(
        n18886) );
  AOI22_X1 U10767 ( .A1(n18300), .A2(n839), .B1(net767235), .B2(net741388), 
        .ZN(n18879) );
  AOI22_X1 U10768 ( .A1(net767167), .A2(n838), .B1(n18326), .B2(net741389), 
        .ZN(n18887) );
  AOI22_X1 U10770 ( .A1(n18330), .A2(n843), .B1(n18331), .B2(n17766), .ZN(
        n18885) );
  INV_X1 U10868 ( .A(n18361), .ZN(n18339) );
  INV_X1 U10869 ( .A(n18369), .ZN(n18338) );
  AOI22_X1 U10756 ( .A1(n18338), .A2(n845), .B1(n18339), .B2(n842), .ZN(n18870) );
  OAI22_X1 U10754 ( .A1(n860), .A2(net767237), .B1(net716477), .B2(net741520), 
        .ZN(n18873) );
  NOR2_X1 U10755 ( .A1(n861), .A2(net767232), .ZN(n18872) );
  AOI211_X1 U10753 ( .C1(n836), .C2(n18343), .A(n18872), .B(n18873), .ZN(
        n18871) );
  AOI22_X1 U10757 ( .A1(net716461), .A2(n841), .B1(n18347), .B2(n847), .ZN(
        n18869) );
  INV_X1 U10944 ( .A(n18393), .ZN(n18311) );
  INV_X1 U10945 ( .A(n18382), .ZN(n18310) );
  AOI22_X1 U10766 ( .A1(n18310), .A2(n851), .B1(n18311), .B2(n837), .ZN(n18880) );
  INV_X1 U10942 ( .A(n18394), .ZN(n18306) );
  AOI22_X1 U10765 ( .A1(net767239), .A2(net741442), .B1(n18306), .B2(n850), 
        .ZN(n18881) );
  INV_X1 U11065 ( .A(n18388), .ZN(n18307) );
  AOI22_X1 U10764 ( .A1(n18307), .A2(n17769), .B1(net716405), .B2(n17768), 
        .ZN(n18882) );
  NAND2_X1 U10760 ( .A1(n18529), .A2(n840), .ZN(n18878) );
  INV_X1 U10875 ( .A(n18390), .ZN(n18321) );
  AOI22_X1 U10761 ( .A1(net767173), .A2(n846), .B1(n18321), .B2(n848), .ZN(
        n18877) );
  OAI211_X1 U10759 ( .C1(n855), .C2(net518461), .A(n18877), .B(n18878), .ZN(
        n18876) );
  INV_X1 U10879 ( .A(n18373), .ZN(n18316) );
  INV_X1 U10880 ( .A(n18372), .ZN(n18315) );
  OAI22_X1 U10762 ( .A1(n863), .A2(n18315), .B1(n862), .B2(n18316), .ZN(n18875) );
  INV_X1 U10881 ( .A(n18387), .ZN(n18312) );
  AOI211_X1 U10758 ( .C1(n18312), .C2(n849), .A(n18875), .B(n18876), .ZN(
        n18868) );
  NOR3_X1 U15971 ( .A1(net715674), .A2(net717955), .A3(net740706), .ZN(
        net715676) );
  NOR2_X1 U15972 ( .A1(net739743), .A2(net715593), .ZN(net715674) );
  NOR3_X1 U15973 ( .A1(net715691), .A2(net715690), .A3(net749287), .ZN(
        net717955) );
  NAND3_X1 U15974 ( .A1(net715668), .A2(net717843), .A3(net740493), .ZN(
        net715691) );
  NAND3_X1 U15975 ( .A1(net715696), .A2(net742068), .A3(net749363), .ZN(
        net715690) );
  AND2_X1 U15976 ( .A1(net715677), .A2(net742073), .ZN(net749287) );
  AND2_X1 U15977 ( .A1(net739688), .A2(net715676), .ZN(net741847) );
  AND2_X2 U15978 ( .A1(net739688), .A2(net715676), .ZN(net713844) );
  NAND3_X1 U15979 ( .A1(net740183), .A2(net715590), .A3(net750077), .ZN(
        net739743) );
  NAND2_X1 U15980 ( .A1(net715696), .A2(net715663), .ZN(net715593) );
  NOR3_X1 U15981 ( .A1(net715674), .A2(net715673), .A3(s_EX_BOT_MUX), .ZN(
        net715672) );
  AND3_X1 U15982 ( .A1(net740305), .A2(net715688), .A3(net715778), .ZN(
        net740183) );
  AND2_X1 U15983 ( .A1(net718026), .A2(net718093), .ZN(net715590) );
  BUF_X1 U15984 ( .A(net715677), .Z(net750077) );
  INV_X1 U15985 ( .A(net739743), .ZN(net715662) );
  NOR2_X1 U15986 ( .A1(n22613), .A2(n22614), .ZN(net740305) );
  NAND2_X1 U15987 ( .A1(n22618), .A2(n22619), .ZN(n22613) );
  XNOR2_X1 U15988 ( .A(net342960), .B(s_MEMWB_IR[13]), .ZN(n22618) );
  XNOR2_X1 U15989 ( .A(net342852), .B(s_MEMWB_IR[15]), .ZN(n22619) );
  NAND3_X1 U15990 ( .A1(n22616), .A2(n22615), .A3(n22617), .ZN(n22614) );
  XNOR2_X1 U15991 ( .A(net718086), .B(s_MEMWB_IR[11]), .ZN(n22616) );
  XNOR2_X1 U15992 ( .A(net718081), .B(s_MEMWB_IR[14]), .ZN(n22615) );
  XNOR2_X1 U15993 ( .A(net718082), .B(s_MEMWB_IR[12]), .ZN(n22617) );
  NAND4_X1 U15994 ( .A1(net715779), .A2(net715780), .A3(net715781), .A4(
        net715782), .ZN(net715688) );
  AOI22_X1 U15995 ( .A1(net715814), .A2(net740357), .B1(net804492), .B2(
        net740358), .ZN(net715778) );
  NAND2_X1 U15996 ( .A1(net740183), .A2(net742288), .ZN(net715666) );
  XOR2_X1 U15997 ( .A(net718138), .B(net718139), .Z(net715814) );
  AND2_X1 U15998 ( .A1(net749815), .A2(s_MEMWB_IR[30]), .ZN(net740357) );
  NAND3_X1 U15999 ( .A1(n22620), .A2(s_MEMWB_IR[28]), .A3(s_MEMWB_IR[27]), 
        .ZN(net804492) );
  XNOR2_X1 U16000 ( .A(net718111), .B(net718098), .ZN(n22620) );
  AOI21_X1 U16001 ( .B1(net745723), .B2(net718138), .A(n18047), .ZN(net740358)
         );
  INV_X1 U16002 ( .A(net715778), .ZN(net720499) );
  NAND3_X1 U16003 ( .A1(n22620), .A2(s_MEMWB_IR[28]), .A3(s_MEMWB_IR[27]), 
        .ZN(net812287) );
  AND2_X1 U16004 ( .A1(s_EX_BOT_MUX), .A2(net741280), .ZN(net740639) );
  AND2_X1 U16005 ( .A1(net740706), .A2(n18051), .ZN(net725586) );
  OR2_X1 U16006 ( .A1(net715593), .A2(n4344), .ZN(net750079) );
  OR2_X1 U16007 ( .A1(net715592), .A2(net715593), .ZN(net725577) );
  NAND4_X1 U16008 ( .A1(net715668), .A2(net715669), .A3(net715590), .A4(
        net715591), .ZN(net740075) );
  NAND4_X1 U16009 ( .A1(net715590), .A2(net715771), .A3(net715772), .A4(
        net749843), .ZN(net715747) );
  NAND3_X1 U16010 ( .A1(net720498), .A2(net750077), .A3(net742288), .ZN(
        net720497) );
  NOR3_X1 U16011 ( .A1(net720499), .A2(net715688), .A3(net715774), .ZN(
        net720498) );
  AOI22_X1 U16012 ( .A1(net715814), .A2(net740357), .B1(net740358), .B2(
        net812287), .ZN(net742073) );
  INV_X1 U16013 ( .A(net715814), .ZN(net715810) );
  NAND2_X1 U16014 ( .A1(s_MEMWB_IR[28]), .A2(s_MEMWB_IR[29]), .ZN(net715706)
         );
  NAND2_X1 U16015 ( .A1(net718138), .A2(net749529), .ZN(net715707) );
  INV_X1 U16016 ( .A(net718139), .ZN(net745725) );
  INV_X1 U16017 ( .A(s_MEMWB_IR[30]), .ZN(net739296) );
  OAI21_X1 U16018 ( .B1(net718111), .B2(s_MEMWB_IR[27]), .A(net742371), .ZN(
        n22612) );
  NOR2_X1 U16019 ( .A1(net745725), .A2(s_MEMWB_IR[29]), .ZN(net745723) );
  CLKBUF_X1 U16020 ( .A(s_MEMWB_IR[29]), .Z(net749815) );
  CLKBUF_X1 U16021 ( .A(net718098), .Z(net742371) );
  INV_X1 U16022 ( .A(net715661), .ZN(net715696) );
  AOI21_X1 U16023 ( .B1(net742011), .B2(net780579), .A(net717926), .ZN(
        net715663) );
  OAI211_X1 U16024 ( .C1(net742047), .C2(net749987), .A(net715795), .B(
        net715796), .ZN(net718026) );
  AOI22_X1 U16025 ( .A1(net750145), .A2(net89524), .B1(net715769), .B2(
        net741339), .ZN(net718093) );
  NAND2_X1 U16026 ( .A1(net715834), .A2(net715705), .ZN(net715677) );
  NOR2_X1 U16027 ( .A1(net715783), .A2(net715784), .ZN(net715779) );
  XNOR2_X1 U16028 ( .A(net366410), .B(s_MEMWB_IR[14]), .ZN(net715780) );
  XNOR2_X1 U16029 ( .A(net342961), .B(s_MEMWB_IR[13]), .ZN(net715781) );
  XNOR2_X1 U16030 ( .A(net342954), .B(s_MEMWB_IR[12]), .ZN(net715782) );
  NOR3_X1 U16031 ( .A1(net715691), .A2(net715690), .A3(net749287), .ZN(
        net715673) );
  CLKBUF_X1 U16032 ( .A(net715696), .Z(net755255) );
  INV_X1 U16033 ( .A(net715696), .ZN(net718033) );
  NAND2_X1 U16034 ( .A1(net715751), .A2(net715663), .ZN(net715746) );
  BUF_X1 U16035 ( .A(net718026), .Z(net749363) );
  AND2_X1 U16036 ( .A1(net786871), .A2(net718026), .ZN(net742288) );
  INV_X1 U16037 ( .A(net715677), .ZN(net715771) );
  NAND2_X1 U16038 ( .A1(net715677), .A2(net742073), .ZN(net715591) );
  NOR3_X1 U16039 ( .A1(net715810), .A2(n22612), .A3(n18047), .ZN(net715695) );
  NOR3_X1 U16040 ( .A1(net715810), .A2(n22612), .A3(n18047), .ZN(net755063) );
  AND2_X1 U16041 ( .A1(n18047), .A2(net739296), .ZN(net715705) );
  INV_X1 U16042 ( .A(net713680), .ZN(net717509) );
  NAND2_X1 U16043 ( .A1(net724878), .A2(net724877), .ZN(net713680) );
  NAND2_X1 U16044 ( .A1(net717509), .A2(net755214), .ZN(net752497) );
  INV_X1 U16045 ( .A(net717509), .ZN(net717511) );
  NOR2_X1 U16046 ( .A1(n22621), .A2(n22622), .ZN(net724878) );
  OR2_X1 U16047 ( .A1(net741960), .A2(n4385), .ZN(net724877) );
  INV_X1 U16048 ( .A(net713680), .ZN(net750122) );
  AND2_X2 U16049 ( .A1(net713680), .A2(net732423), .ZN(net714248) );
  OAI211_X1 U16050 ( .C1(net718360), .C2(net740649), .A(n22624), .B(n22623), 
        .ZN(n22621) );
  INV_X1 U16051 ( .A(net713847), .ZN(net718360) );
  NAND2_X1 U16052 ( .A1(net741847), .A2(net717454), .ZN(n22624) );
  NAND2_X1 U16053 ( .A1(net717517), .A2(n18050), .ZN(n22623) );
  AND2_X1 U16054 ( .A1(net715672), .A2(net739688), .ZN(net717517) );
  NOR2_X1 U16055 ( .A1(net717107), .A2(n1700), .ZN(n22622) );
  BUF_X1 U16056 ( .A(net717103), .Z(net717107) );
  NAND2_X1 U16057 ( .A1(net724878), .A2(net724877), .ZN(net749316) );
  NAND2_X1 U16058 ( .A1(net742258), .A2(net718032), .ZN(net739688) );
  INV_X1 U16059 ( .A(net741847), .ZN(net718351) );
  NAND2_X1 U16060 ( .A1(net741847), .A2(n17957), .ZN(net715524) );
  OAI222_X1 U16061 ( .A1(net780582), .A2(net780188), .B1(n1692), .B2(net717105), .C1(net718360), .C2(net741572), .ZN(net741980) );
  INV_X1 U16062 ( .A(net718360), .ZN(net717789) );
  AOI22_X1 U16063 ( .A1(net741608), .A2(net741464), .B1(net712606), .B2(n5707), 
        .ZN(net715892) );
  AOI22_X1 U16064 ( .A1(net755033), .A2(n5707), .B1(net742412), .B2(
        \core_inst/MEMWB_ALUOUT/DFF_2/N3 ), .ZN(net736610) );
  NOR2_X1 U16065 ( .A1(net716311), .A2(n5601), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_2/N3 ) );
  AND2_X1 U16066 ( .A1(net715672), .A2(net739688), .ZN(net762579) );
  NAND2_X1 U16067 ( .A1(net715647), .A2(net717742), .ZN(net741960) );
  AND3_X1 U16068 ( .A1(net742257), .A2(net765400), .A3(net750053), .ZN(
        net713847) );
  NAND2_X1 U16069 ( .A1(net762761), .A2(net715700), .ZN(net742258) );
  AND2_X2 U16070 ( .A1(net755255), .A2(net718092), .ZN(net718032) );
  BUF_X1 U16071 ( .A(net741960), .Z(net741959) );
  BUF_X1 U16072 ( .A(net741960), .Z(net741958) );
  NAND2_X1 U16073 ( .A1(net750031), .A2(net741464), .ZN(net736609) );
  OAI22_X1 U16074 ( .A1(net717107), .A2(n1694), .B1(net714943), .B2(net740661), 
        .ZN(net715221) );
  OAI222_X1 U16075 ( .A1(net718351), .A2(net780188), .B1(net717107), .B2(n1692), .C1(net718361), .C2(net741572), .ZN(net715603) );
  INV_X1 U16076 ( .A(net713847), .ZN(net718361) );
  INV_X1 U16077 ( .A(net717517), .ZN(net738474) );
  NAND2_X1 U16078 ( .A1(net742258), .A2(net718032), .ZN(net717742) );
  NAND3_X1 U16079 ( .A1(net715656), .A2(net742257), .A3(net718032), .ZN(
        net717104) );
  NAND3_X1 U16080 ( .A1(net715656), .A2(net742257), .A3(net718032), .ZN(
        net717103) );
  NOR4_X1 U16081 ( .A1(net712799), .A2(net713453), .A3(net712815), .A4(
        net712452), .ZN(n22625) );
  OAI211_X1 U16082 ( .C1(net714406), .C2(net713751), .A(net714408), .B(
        net714407), .ZN(net712799) );
  OAI211_X1 U16083 ( .C1(net714375), .C2(net713751), .A(net714376), .B(
        net714377), .ZN(net713453) );
  NAND3_X1 U16084 ( .A1(net727827), .A2(net727829), .A3(net727828), .ZN(
        net712815) );
  OAI211_X1 U16085 ( .C1(net714360), .C2(net767203), .A(net714361), .B(
        net714362), .ZN(net712452) );
  NAND3_X1 U16086 ( .A1(net740705), .A2(net713062), .A3(n22625), .ZN(net714332) );
  NOR4_X1 U16087 ( .A1(n22632), .A2(n22631), .A3(n22633), .A4(n22634), .ZN(
        net714360) );
  OAI222_X1 U16088 ( .A1(net717055), .A2(net755238), .B1(net717075), .B2(
        net749525), .C1(net728314), .C2(net749823), .ZN(n22632) );
  CLKBUF_X3 U16089 ( .A(net713866), .Z(net717055) );
  CLKBUF_X3 U16090 ( .A(net714251), .Z(net755238) );
  CLKBUF_X3 U16091 ( .A(net712470), .Z(net717075) );
  CLKBUF_X1 U16092 ( .A(net767335), .Z(net749525) );
  NAND2_X2 U16093 ( .A1(net717463), .A2(net713733), .ZN(net728314) );
  INV_X1 U16094 ( .A(net749820), .ZN(net749823) );
  OAI222_X1 U16095 ( .A1(net713907), .A2(net713681), .B1(net718406), .B2(
        net749260), .C1(net750278), .C2(net767207), .ZN(n22631) );
  NAND2_X2 U16096 ( .A1(net749372), .A2(net715284), .ZN(net713907) );
  INV_X1 U16097 ( .A(net755610), .ZN(net713681) );
  BUF_X1 U16098 ( .A(net713853), .Z(net718406) );
  NAND2_X1 U16099 ( .A1(net767352), .A2(net740674), .ZN(net749260) );
  NAND2_X1 U16100 ( .A1(net755048), .A2(net742248), .ZN(net750278) );
  INV_X1 U16101 ( .A(net714194), .ZN(net767207) );
  OAI22_X1 U16102 ( .A1(net750274), .A2(net717053), .B1(net713851), .B2(
        net742271), .ZN(n22633) );
  INV_X1 U16103 ( .A(net713687), .ZN(net750274) );
  BUF_X2 U16104 ( .A(net712893), .Z(net717053) );
  OR2_X1 U16105 ( .A1(net750203), .A2(net737907), .ZN(net713851) );
  INV_X1 U16106 ( .A(net713683), .ZN(net742271) );
  OAI22_X1 U16107 ( .A1(net717059), .A2(net750093), .B1(net717875), .B2(
        net748275), .ZN(n22634) );
  BUF_X2 U16108 ( .A(net713864), .Z(net717059) );
  INV_X1 U16109 ( .A(net749832), .ZN(net750093) );
  CLKBUF_X3 U16110 ( .A(net750228), .Z(net717875) );
  INV_X1 U16111 ( .A(net737713), .ZN(net748275) );
  INV_X1 U16112 ( .A(net713775), .ZN(net767203) );
  NOR2_X1 U16113 ( .A1(n22626), .A2(n22627), .ZN(net714361) );
  AND2_X1 U16114 ( .A1(n22638), .A2(net714876), .ZN(n22626) );
  AND4_X1 U16115 ( .A1(net714873), .A2(net714877), .A3(net714275), .A4(
        net753553), .ZN(n22638) );
  NAND2_X1 U16116 ( .A1(net763705), .A2(net714476), .ZN(net714873) );
  NAND2_X1 U16117 ( .A1(net749886), .A2(net750238), .ZN(net714877) );
  AND2_X2 U16118 ( .A1(net713733), .A2(net767221), .ZN(net714275) );
  NAND2_X1 U16119 ( .A1(net717464), .A2(net713753), .ZN(net753553) );
  AOI21_X1 U16120 ( .B1(net750158), .B2(net742507), .A(net786066), .ZN(
        net714876) );
  OAI21_X1 U16121 ( .B1(n22641), .B2(net767210), .A(n22628), .ZN(n22627) );
  NAND4_X1 U16122 ( .A1(n22636), .A2(n22635), .A3(n22637), .A4(net714965), 
        .ZN(n22641) );
  AOI22_X1 U16123 ( .A1(net713773), .A2(net714967), .B1(n22642), .B2(net750019), .ZN(n22636) );
  AOI22_X1 U16124 ( .A1(net714874), .A2(net718355), .B1(net750159), .B2(
        net718391), .ZN(n22635) );
  AOI22_X1 U16125 ( .A1(net717464), .A2(net749306), .B1(net742157), .B2(
        net750251), .ZN(n22637) );
  NAND2_X1 U16126 ( .A1(net714476), .A2(net718025), .ZN(net714965) );
  INV_X1 U16127 ( .A(net714309), .ZN(net767210) );
  MUX2_X1 U16128 ( .A(n22629), .B(n22630), .S(net717875), .Z(n22628) );
  MUX2_X1 U16129 ( .A(net713726), .B(net713738), .S(net755090), .Z(n22629) );
  NAND2_X1 U16130 ( .A1(net715584), .A2(net716231), .ZN(net713726) );
  NAND2_X1 U16131 ( .A1(net715584), .A2(net741282), .ZN(net713738) );
  AND2_X1 U16132 ( .A1(net780568), .A2(net715175), .ZN(net755090) );
  MUX2_X1 U16133 ( .A(net713728), .B(net717087), .S(net755090), .Z(n22630) );
  NAND2_X2 U16134 ( .A1(net715584), .A2(net741531), .ZN(net713728) );
  NAND2_X1 U16135 ( .A1(net715584), .A2(net741603), .ZN(net717087) );
  INV_X1 U16136 ( .A(net795965), .ZN(net714362) );
  OAI33_X1 U16137 ( .A1(n22640), .A2(net715015), .A3(net795964), .B1(net715236), .B2(net715235), .B3(net714267), .ZN(net795965) );
  NAND4_X1 U16138 ( .A1(net731685), .A2(net715018), .A3(net715019), .A4(
        net715020), .ZN(n22640) );
  AND2_X1 U16139 ( .A1(net715014), .A2(net715021), .ZN(net731685) );
  NAND2_X1 U16140 ( .A1(net749317), .A2(net717875), .ZN(net715018) );
  NAND2_X1 U16141 ( .A1(net714874), .A2(net755241), .ZN(net715019) );
  NAND2_X1 U16142 ( .A1(net750159), .A2(net713614), .ZN(net715020) );
  NAND2_X1 U16143 ( .A1(net714965), .A2(net715232), .ZN(net715015) );
  INV_X1 U16144 ( .A(net714306), .ZN(net795964) );
  AND2_X1 U16145 ( .A1(net715313), .A2(net713863), .ZN(net714306) );
  OR3_X1 U16146 ( .A1(net717778), .A2(net717779), .A3(net717780), .ZN(
        net715236) );
  NAND3_X1 U16147 ( .A1(n22643), .A2(net781609), .A3(net714965), .ZN(net715235) );
  NAND2_X1 U16148 ( .A1(net715284), .A2(net713863), .ZN(net714267) );
  CLKBUF_X1 U16149 ( .A(net712452), .Z(net742100) );
  MUX2_X2 U16150 ( .A(n478), .B(net714078), .S(net716237), .Z(net713773) );
  INV_X1 U16151 ( .A(net715242), .ZN(net714967) );
  BUF_X1 U16152 ( .A(n22639), .Z(n22642) );
  MUX2_X2 U16153 ( .A(net762727), .B(n13805), .S(net741686), .Z(net750019) );
  NAND4_X1 U16154 ( .A1(n22636), .A2(n22635), .A3(n22637), .A4(net714965), 
        .ZN(net714344) );
  NOR2_X1 U16155 ( .A1(net752497), .A2(net742243), .ZN(n22639) );
  AOI22_X1 U16156 ( .A1(n22642), .A2(net742315), .B1(net714967), .B2(net748274), .ZN(n22643) );
  INV_X1 U16157 ( .A(n22642), .ZN(net749902) );
  BUF_X2 U16158 ( .A(net755262), .Z(net742243) );
  CLKBUF_X1 U16159 ( .A(n22639), .Z(net749500) );
  OR2_X2 U16160 ( .A1(net715603), .A2(net737941), .ZN(net755214) );
  NOR2_X1 U16161 ( .A1(net742243), .A2(net752497), .ZN(net749886) );
  NOR2_X1 U16162 ( .A1(net752497), .A2(net749697), .ZN(net749372) );
  CLKBUF_X1 U16163 ( .A(net712799), .Z(net742182) );
  CLKBUF_X1 U16164 ( .A(net713453), .Z(net717654) );
  CLKBUF_X1 U16165 ( .A(net712815), .Z(net780551) );
  NAND2_X1 U16166 ( .A1(net714967), .A2(net713868), .ZN(net715241) );
  NAND2_X1 U16167 ( .A1(net714967), .A2(net742087), .ZN(net715232) );
  NOR4_X1 U16168 ( .A1(net714431), .A2(net714433), .A3(net714432), .A4(
        net714434), .ZN(net714406) );
  INV_X1 U16169 ( .A(net713863), .ZN(net713751) );
  MUX2_X1 U16170 ( .A(net714409), .B(net714410), .S(net718380), .Z(net714408)
         );
  NOR3_X1 U16171 ( .A1(net714415), .A2(net714414), .A3(net714413), .ZN(
        net714407) );
  NOR4_X1 U16172 ( .A1(net714386), .A2(net714387), .A3(net714389), .A4(
        net714388), .ZN(net714375) );
  NOR2_X1 U16173 ( .A1(net714379), .A2(net714380), .ZN(net714376) );
  NAND2_X1 U16174 ( .A1(net714378), .A2(net739078), .ZN(net714377) );
  AOI22_X1 U16175 ( .A1(net713978), .A2(net713785), .B1(net713979), .B2(
        net767211), .ZN(net727827) );
  NOR2_X1 U16176 ( .A1(net727830), .A2(net727831), .ZN(net727829) );
  OAI21_X1 U16177 ( .B1(net727833), .B2(net727834), .A(net767221), .ZN(
        net727828) );
  NOR3_X4 U16178 ( .A1(net366451), .A2(net366531), .A3(net366479), .ZN(
        net713775) );
  AND2_X1 U16179 ( .A1(net713740), .A2(net713863), .ZN(net714309) );
  BUF_X1 U16180 ( .A(net731344), .Z(net714874) );
  CLKBUF_X1 U16181 ( .A(net755216), .Z(net718355) );
  AND2_X2 U16182 ( .A1(net762604), .A2(net747343), .ZN(net750159) );
  CLKBUF_X3 U16183 ( .A(net713777), .Z(net718391) );
  INV_X1 U16184 ( .A(net717461), .ZN(net717464) );
  MUX2_X2 U16185 ( .A(n1182), .B(net749308), .S(net787512), .Z(net749306) );
  MUX2_X2 U16186 ( .A(n1064), .B(net714077), .S(net787518), .Z(net742157) );
  NOR2_X1 U16187 ( .A1(net765428), .A2(net742243), .ZN(net750251) );
  OR2_X2 U16188 ( .A1(net718349), .A2(net741282), .ZN(net714476) );
  INV_X1 U16189 ( .A(net749465), .ZN(net718025) );
  NOR2_X1 U16190 ( .A1(net715575), .A2(net715576), .ZN(net714078) );
  INV_X2 U16191 ( .A(net741686), .ZN(net716237) );
  NAND2_X1 U16192 ( .A1(net714248), .A2(net742242), .ZN(net715242) );
  NOR2_X1 U16193 ( .A1(net765677), .A2(net747437), .ZN(net762727) );
  OR2_X1 U16194 ( .A1(net715586), .A2(net715528), .ZN(net755262) );
  OAI22_X1 U16195 ( .A1(net737101), .A2(n4352), .B1(net738474), .B2(net741306), 
        .ZN(net737941) );
  AND2_X1 U16196 ( .A1(net714876), .A2(net749427), .ZN(net714657) );
  AND2_X1 U16197 ( .A1(net714876), .A2(net767208), .ZN(net733229) );
  AOI222_X1 U16198 ( .A1(net742157), .A2(net750159), .B1(net742247), .B2(
        net749525), .C1(net749489), .C2(net767207), .ZN(net715555) );
  NAND2_X1 U16199 ( .A1(net750159), .A2(net718380), .ZN(net715027) );
  INV_X1 U16200 ( .A(net750251), .ZN(net755683) );
  INV_X1 U16201 ( .A(net718025), .ZN(net782764) );
  NAND2_X1 U16202 ( .A1(net713679), .A2(net718025), .ZN(net715333) );
  MUX2_X2 U16203 ( .A(n478), .B(net714078), .S(net787518), .Z(net718349) );
  CLKBUF_X1 U16204 ( .A(net714078), .Z(net762762) );
  NOR2_X1 U16205 ( .A1(net715242), .A2(net714559), .ZN(net784601) );
  BUF_X1 U16206 ( .A(net715242), .Z(net762729) );
  MUX2_X1 U16207 ( .A(net714076), .B(n13805), .S(net741686), .Z(net713627) );
  INV_X1 U16208 ( .A(net741726), .ZN(net787514) );
  BUF_X1 U16209 ( .A(net741726), .Z(net787512) );
  INV_X1 U16210 ( .A(net741726), .ZN(net787516) );
  MUX2_X1 U16211 ( .A(n367), .B(net742224), .S(net741726), .Z(net713709) );
  BUF_X2 U16212 ( .A(net755262), .Z(net742242) );
  BUF_X1 U16213 ( .A(net755262), .Z(net749698) );
  CLKBUF_X1 U16214 ( .A(net715603), .Z(net786852) );
  NOR2_X1 U16215 ( .A1(net737937), .A2(net715603), .ZN(net749375) );
  NOR2_X1 U16216 ( .A1(net741980), .A2(net737941), .ZN(net732423) );
  OAI21_X1 U16217 ( .B1(net804645), .B2(n22645), .A(n22646), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_20/N3 ) );
  INV_X1 U16218 ( .A(net716387), .ZN(net804645) );
  OAI21_X1 U16219 ( .B1(n22647), .B2(n22648), .A(net717052), .ZN(n22645) );
  NAND4_X1 U16220 ( .A1(n18868), .A2(n22663), .A3(n18869), .A4(n22651), .ZN(
        n22647) );
  NAND2_X1 U16221 ( .A1(net715842), .A2(n19255), .ZN(net518461) );
  INV_X1 U16222 ( .A(n18400), .ZN(net767173) );
  INV_X1 U16223 ( .A(n18318), .ZN(n18529) );
  AND3_X1 U16224 ( .A1(n18882), .A2(n18881), .A3(n18880), .ZN(n22663) );
  INV_X2 U16225 ( .A(net741549), .ZN(net716405) );
  INV_X2 U16226 ( .A(net741541), .ZN(net767239) );
  INV_X2 U16227 ( .A(n18346), .ZN(net716461) );
  NOR2_X2 U16228 ( .A1(net708964), .A2(n19245), .ZN(n18347) );
  AND2_X1 U16229 ( .A1(n18871), .A2(n18870), .ZN(n22651) );
  NOR2_X2 U16230 ( .A1(n19262), .A2(n19248), .ZN(n18343) );
  INV_X2 U16231 ( .A(net716491), .ZN(net767232) );
  INV_X2 U16232 ( .A(net741532), .ZN(net767237) );
  INV_X2 U16233 ( .A(net741539), .ZN(net716477) );
  NAND4_X1 U16234 ( .A1(n22662), .A2(n18887), .A3(n18879), .A4(n18886), .ZN(
        n22648) );
  AND3_X1 U16235 ( .A1(n18885), .A2(n22649), .A3(n22650), .ZN(n22662) );
  INV_X2 U16236 ( .A(n18362), .ZN(n18330) );
  INV_X1 U16237 ( .A(n18363), .ZN(n18331) );
  OR2_X1 U16238 ( .A1(n18332), .A2(n858), .ZN(n22649) );
  NAND2_X2 U16239 ( .A1(n19255), .A2(n19242), .ZN(n18332) );
  NAND2_X1 U16240 ( .A1(n18398), .A2(net741397), .ZN(n22650) );
  NOR2_X1 U16241 ( .A1(n19248), .A2(n19261), .ZN(n18398) );
  BUF_X2 U16242 ( .A(n18325), .Z(net767167) );
  NOR2_X2 U16243 ( .A1(n19248), .A2(n19245), .ZN(n18326) );
  INV_X1 U16244 ( .A(n18395), .ZN(n18300) );
  INV_X2 U16245 ( .A(net741544), .ZN(net767235) );
  NOR2_X2 U16246 ( .A1(n19262), .A2(n19246), .ZN(n18328) );
  AND2_X1 U16247 ( .A1(net713412), .A2(net713414), .ZN(net717052) );
  NAND2_X1 U16248 ( .A1(net716255), .A2(n22666), .ZN(n22646) );
  INV_X1 U16249 ( .A(net795260), .ZN(net716255) );
  AND2_X1 U16250 ( .A1(net717049), .A2(net712946), .ZN(n22666) );
  AND2_X1 U16251 ( .A1(net713412), .A2(net713413), .ZN(net717049) );
  INV_X1 U16252 ( .A(net717157), .ZN(net712946) );
  BUF_X1 U16253 ( .A(net717950), .Z(net795260) );
  AND2_X1 U16254 ( .A1(n22653), .A2(net760672), .ZN(net717950) );
  INV_X1 U16255 ( .A(net795260), .ZN(net716259) );
  INV_X1 U16256 ( .A(net795260), .ZN(net741999) );
  OAI21_X1 U16257 ( .B1(net714030), .B2(net714031), .A(net713490), .ZN(n22653)
         );
  OAI22_X1 U16258 ( .A1(net713488), .A2(net760673), .B1(net713490), .B2(
        net740645), .ZN(net760672) );
  NAND3_X1 U16259 ( .A1(net714619), .A2(net714621), .A3(net714620), .ZN(
        net714030) );
  NAND4_X1 U16260 ( .A1(net714085), .A2(net714086), .A3(net780225), .A4(
        net714087), .ZN(net714031) );
  XNOR2_X1 U16261 ( .A(net714032), .B(s_EX_BRANCH_TYPE), .ZN(net713490) );
  CLKBUF_X1 U16262 ( .A(n22653), .Z(net780532) );
  NOR3_X1 U16263 ( .A1(n22657), .A2(net714332), .A3(net714330), .ZN(net714085)
         );
  NAND4_X1 U16264 ( .A1(net712888), .A2(n22659), .A3(net713461), .A4(net713455), .ZN(n22657) );
  OAI211_X1 U16265 ( .C1(net714529), .C2(net714530), .A(net714532), .B(
        net714531), .ZN(net712888) );
  NOR2_X1 U16266 ( .A1(net713208), .A2(n22644), .ZN(n22659) );
  NAND4_X1 U16267 ( .A1(net714506), .A2(net714508), .A3(net714507), .A4(
        net746315), .ZN(net713208) );
  NAND4_X1 U16268 ( .A1(net714486), .A2(net714487), .A3(net714488), .A4(
        net714489), .ZN(n22644) );
  NOR2_X1 U16269 ( .A1(net714501), .A2(net714502), .ZN(net714486) );
  AOI22_X1 U16270 ( .A1(net713873), .A2(net713779), .B1(net713870), .B2(
        net713785), .ZN(net714487) );
  MUX2_X1 U16271 ( .A(net714492), .B(net714493), .S(net714494), .Z(net714488)
         );
  OAI21_X1 U16272 ( .B1(net714490), .B2(net714491), .A(net713863), .ZN(
        net714489) );
  OAI211_X1 U16273 ( .C1(net714463), .C2(net714464), .A(net714465), .B(
        net714466), .ZN(net713461) );
  NAND3_X1 U16274 ( .A1(net729531), .A2(net725022), .A3(net729530), .ZN(
        net713455) );
  AND2_X1 U16275 ( .A1(net712559), .A2(n22658), .ZN(net740705) );
  OAI211_X1 U16276 ( .C1(net738840), .C2(net724910), .A(net738839), .B(
        net717091), .ZN(net712559) );
  NAND3_X1 U16277 ( .A1(net733097), .A2(net717091), .A3(net713463), .ZN(n22658) );
  OAI21_X1 U16278 ( .B1(net755783), .B2(net714337), .A(net713469), .ZN(
        net733097) );
  BUF_X2 U16279 ( .A(net712459), .Z(net717091) );
  INV_X1 U16280 ( .A(net714335), .ZN(net713463) );
  NOR4_X1 U16281 ( .A1(net714339), .A2(net714340), .A3(net714341), .A4(
        net714342), .ZN(net713062) );
  OAI211_X1 U16282 ( .C1(net767210), .C2(net714354), .A(net714355), .B(
        net714356), .ZN(net714339) );
  AOI21_X1 U16283 ( .B1(net714346), .B2(net714347), .A(net767203), .ZN(
        net714340) );
  NOR2_X1 U16284 ( .A1(net713692), .A2(net713738), .ZN(net714341) );
  OAI21_X1 U16285 ( .B1(net714344), .B2(net767209), .A(net733227), .ZN(
        net714342) );
  OAI21_X1 U16286 ( .B1(net713067), .B2(net727306), .A(net713068), .ZN(
        net714330) );
  NOR2_X1 U16287 ( .A1(n22654), .A2(n22660), .ZN(net714086) );
  NAND3_X1 U16288 ( .A1(n22655), .A2(n22652), .A3(n22656), .ZN(n22654) );
  NOR2_X1 U16289 ( .A1(net731393), .A2(net731713), .ZN(n22655) );
  NAND2_X1 U16290 ( .A1(net717684), .A2(net749219), .ZN(net731393) );
  AOI21_X1 U16291 ( .B1(net733282), .B2(net733283), .A(net713154), .ZN(
        net731713) );
  NAND2_X1 U16292 ( .A1(net734282), .A2(net717091), .ZN(n22652) );
  XNOR2_X1 U16293 ( .A(net783466), .B(net783467), .ZN(net734282) );
  NOR3_X1 U16294 ( .A1(net712931), .A2(net712856), .A3(n22661), .ZN(n22656) );
  NAND4_X1 U16295 ( .A1(net714172), .A2(net714174), .A3(net714173), .A4(
        net714175), .ZN(net712931) );
  NAND3_X1 U16296 ( .A1(net778055), .A2(net778056), .A3(net778057), .ZN(
        net712856) );
  NAND2_X1 U16297 ( .A1(n22664), .A2(net758544), .ZN(n22661) );
  AND2_X1 U16298 ( .A1(net714239), .A2(n22665), .ZN(n22664) );
  AOI21_X1 U16299 ( .B1(net714240), .B2(net767211), .A(net714241), .ZN(
        net714239) );
  INV_X1 U16300 ( .A(net712857), .ZN(n22665) );
  NOR2_X1 U16301 ( .A1(net714227), .A2(net714228), .ZN(net712857) );
  NAND2_X1 U16302 ( .A1(net729177), .A2(net729185), .ZN(net758544) );
  OR2_X1 U16303 ( .A1(net737706), .A2(net738517), .ZN(n22660) );
  NOR2_X1 U16304 ( .A1(net714140), .A2(net737707), .ZN(net737706) );
  AOI21_X1 U16305 ( .B1(net745867), .B2(net745868), .A(net713154), .ZN(
        net738517) );
  NAND2_X1 U16306 ( .A1(net729283), .A2(net729282), .ZN(net780225) );
  NAND3_X1 U16307 ( .A1(net713449), .A2(net717091), .A3(net713450), .ZN(
        net714087) );
  NAND2_X1 U16308 ( .A1(net714106), .A2(net749533), .ZN(net713449) );
  INV_X1 U16309 ( .A(net714105), .ZN(net713450) );
  OAI21_X1 U16310 ( .B1(net714030), .B2(net714031), .A(net713490), .ZN(
        net765379) );
  NOR2_X1 U16311 ( .A1(net804645), .A2(net873523), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_10/N3 ) );
  NOR2_X1 U16312 ( .A1(net804645), .A2(net780186), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_21/N3 ) );
  AND2_X1 U16313 ( .A1(net765379), .A2(net760672), .ZN(net765340) );
  OAI22_X1 U16314 ( .A1(net755203), .A2(net755094), .B1(net713490), .B2(
        net740645), .ZN(net755005) );
  CLKBUF_X1 U16315 ( .A(net780225), .Z(net796204) );
  CLKBUF_X1 U16316 ( .A(net714330), .Z(net749292) );
  BUF_X1 U16317 ( .A(n15091), .Z(net716387) );
  NAND3_X1 U16318 ( .A1(net713757), .A2(net713756), .A3(net713755), .ZN(
        net713488) );
  AOI22_X1 U16319 ( .A1(net713492), .A2(net712966), .B1(net713493), .B2(
        net713494), .ZN(net760673) );
  NOR3_X1 U16320 ( .A1(net714909), .A2(net714910), .A3(net714911), .ZN(
        net714619) );
  NOR2_X1 U16321 ( .A1(net714622), .A2(net713442), .ZN(net714621) );
  NOR3_X1 U16322 ( .A1(net714732), .A2(net712445), .A3(net740704), .ZN(
        net714620) );
  NOR2_X1 U16323 ( .A1(net714033), .A2(net714034), .ZN(net714032) );
  OAI21_X1 U16324 ( .B1(net714096), .B2(net749533), .A(net729284), .ZN(
        net729283) );
  NAND3_X1 U16325 ( .A1(net729291), .A2(net729292), .A3(net749454), .ZN(
        net729282) );
  AOI21_X1 U16326 ( .B1(net720369), .B2(net720368), .A(net720370), .ZN(
        net713067) );
  NAND2_X1 U16327 ( .A1(net725126), .A2(net725127), .ZN(net727306) );
  NOR3_X1 U16328 ( .A1(net714552), .A2(net714553), .A3(net740679), .ZN(
        net713068) );
  AND2_X1 U16329 ( .A1(net717048), .A2(net712946), .ZN(net712945) );
  CLKBUF_X1 U16330 ( .A(net713488), .Z(net755203) );
  NAND3_X1 U16331 ( .A1(net726729), .A2(s_EX_IS_BRANCH), .A3(net713074), .ZN(
        net713758) );
  MUX2_X1 U16332 ( .A(net713448), .B(net713449), .S(net713450), .Z(net713446)
         );
  CLKBUF_X1 U16333 ( .A(net712888), .Z(net780537) );
  CLKBUF_X1 U16334 ( .A(net713461), .Z(net780599) );
  OAI21_X1 U16335 ( .B1(net780337), .B2(net717696), .A(net713455), .ZN(
        net780338) );
  INV_X1 U16336 ( .A(net712559), .ZN(net742198) );
  OR4_X1 U16337 ( .A1(net714340), .A2(net714339), .A3(net714342), .A4(
        net714341), .ZN(net780214) );
  MUX2_X1 U16338 ( .A(n26078), .B(n1182), .S(net787516), .Z(net765546) );
  INV_X2 U16339 ( .A(net787516), .ZN(net787518) );
  CLKBUF_X1 U16340 ( .A(n25853), .Z(n22667) );
  INV_X1 U16341 ( .A(net762579), .ZN(net767340) );
  INV_X1 U16342 ( .A(n22669), .ZN(n22675) );
  OR2_X1 U16344 ( .A1(n26637), .A2(n26630), .ZN(n22670) );
  OR2_X1 U16345 ( .A1(n26637), .A2(n26447), .ZN(n22671) );
  OR2_X2 U16346 ( .A1(net796126), .A2(net786852), .ZN(n22673) );
  CLKBUF_X1 U16347 ( .A(net715445), .Z(net749408) );
  AND2_X1 U16348 ( .A1(net717050), .A2(n26467), .ZN(n22678) );
  AND2_X1 U16349 ( .A1(net717050), .A2(n26661), .ZN(n22679) );
  AND2_X1 U16350 ( .A1(n25665), .A2(n26299), .ZN(n22680) );
  AND2_X1 U16351 ( .A1(net712397), .A2(n26400), .ZN(n22681) );
  OR2_X1 U16352 ( .A1(n23138), .A2(n23139), .ZN(n22682) );
  INV_X1 U16353 ( .A(n24547), .ZN(n22980) );
  AND2_X1 U16354 ( .A1(n18136), .A2(n25336), .ZN(n22683) );
  AND2_X1 U16355 ( .A1(n26599), .A2(n25664), .ZN(n22684) );
  AND2_X1 U16356 ( .A1(net718074), .A2(s_IFID_IR[16]), .ZN(n22685) );
  NAND2_X1 U16357 ( .A1(net717050), .A2(n26631), .ZN(n22689) );
  NAND2_X1 U16358 ( .A1(n25665), .A2(n26631), .ZN(n22690) );
  NAND2_X1 U16359 ( .A1(net717048), .A2(n26448), .ZN(n22691) );
  OAI21_X1 U16361 ( .B1(net712367), .B2(net716263), .A(n22693), .ZN(net521855)
         );
  AOI21_X1 U16362 ( .B1(net717091), .B2(net780294), .A(net780295), .ZN(
        net712367) );
  INV_X1 U16363 ( .A(net716339), .ZN(net716263) );
  NAND2_X1 U16364 ( .A1(net716251), .A2(n22694), .ZN(n22693) );
  INV_X1 U16365 ( .A(net717967), .ZN(net716251) );
  INV_X1 U16366 ( .A(n22695), .ZN(n22694) );
  OAI21_X1 U16367 ( .B1(net785319), .B2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [28]), .A(net712847), .ZN(n22695) );
  NOR3_X1 U16368 ( .A1(net712838), .A2(n6402), .A3(net780340), .ZN(net785319)
         );
  NAND2_X1 U16369 ( .A1(net712886), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [28]), .ZN(net712847) );
  INV_X1 U16370 ( .A(n22693), .ZN(net812861) );
  CLKBUF_X2 U16371 ( .A(net717950), .Z(net717967) );
  NAND2_X1 U16372 ( .A1(net716251), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [1]), .ZN(net712391) );
  NAND2_X1 U16373 ( .A1(net716251), .A2(s_IFID_IR[21]), .ZN(net712384) );
  NAND2_X1 U16374 ( .A1(net716251), .A2(n18136), .ZN(net812773) );
  NOR2_X1 U16375 ( .A1(net785270), .A2(net712367), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_28/N3 ) );
  OAI21_X1 U16376 ( .B1(net713463), .B2(net780291), .A(net780293), .ZN(
        net780294) );
  INV_X1 U16377 ( .A(net780599), .ZN(net780295) );
  CLKBUF_X3 U16378 ( .A(net765340), .Z(net716339) );
  CLKBUF_X3 U16379 ( .A(net795568), .Z(net796232) );
  CLKBUF_X1 U16380 ( .A(n25872), .Z(n22696) );
  CLKBUF_X3 U16381 ( .A(net716337), .Z(net796143) );
  INV_X1 U16382 ( .A(n26744), .ZN(n22704) );
  OAI21_X1 U16383 ( .B1(net716263), .B2(net712366), .A(n22697), .ZN(n16388) );
  NOR2_X1 U16384 ( .A1(net717654), .A2(net780338), .ZN(net712366) );
  NAND2_X1 U16385 ( .A1(net796255), .A2(net713451), .ZN(n22697) );
  INV_X1 U16386 ( .A(net716337), .ZN(net796255) );
  AOI21_X1 U16387 ( .B1(n6512), .B2(net713441), .A(net712795), .ZN(net713451)
         );
  CLKBUF_X2 U16388 ( .A(net717950), .Z(net716337) );
  NOR2_X1 U16389 ( .A1(net716313), .A2(net712366), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_19/N3 ) );
  AND2_X1 U16390 ( .A1(net785255), .A2(net713451), .ZN(net780182) );
  NAND2_X1 U16391 ( .A1(net712922), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [18]), .ZN(net713441) );
  NOR2_X2 U16392 ( .A1(net713441), .A2(n6512), .ZN(net712795) );
  OAI21_X1 U16393 ( .B1(net712922), .B2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [18]), .A(net713441), .ZN(net713439) );
  OR2_X1 U16394 ( .A1(net717967), .A2(n23536), .ZN(n22874) );
  NAND2_X1 U16395 ( .A1(net716259), .A2(n22678), .ZN(n24436) );
  BUF_X1 U16396 ( .A(net717720), .Z(net718340) );
  OR2_X1 U16397 ( .A1(net796271), .A2(net741237), .ZN(n13343) );
  AND2_X1 U16398 ( .A1(net716243), .A2(n22941), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_19/N3 ) );
  NOR2_X1 U16399 ( .A1(net796143), .A2(n22698), .ZN(
        \core_inst/IDEX_NPC/DFF_4/N3 ) );
  NOR2_X1 U16400 ( .A1(net796143), .A2(n24618), .ZN(n22801) );
  NOR2_X1 U16401 ( .A1(net796143), .A2(n22699), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_6/N3 ) );
  NOR2_X1 U16402 ( .A1(net796133), .A2(n22700), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_11/N3 ) );
  INV_X32 U16403 ( .A(n22943), .ZN(n22700) );
  NOR2_X1 U16404 ( .A1(net796232), .A2(n22701), .ZN(
        \core_inst/IDEX_NPC/DFF_28/N3 ) );
  BUF_X1 U16405 ( .A(net717967), .Z(net716331) );
  AND2_X1 U16406 ( .A1(net741999), .A2(s_IFID_IR[24]), .ZN(n22702) );
  AND2_X1 U16407 ( .A1(net760161), .A2(s_IFID_IR[18]), .ZN(n22703) );
  NOR2_X1 U16408 ( .A1(net716313), .A2(n24612), .ZN(
        \core_inst/IDEX_IR/DFF_31/N3 ) );
  NOR2_X1 U16409 ( .A1(net716333), .A2(n22704), .ZN(
        \core_inst/IFID_NPC/DFF_3/N3 ) );
  AND2_X1 U16410 ( .A1(net716257), .A2(net839583), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_1/N3 ) );
  INV_X32 U16411 ( .A(n1501), .ZN(net839583) );
  AND2_X1 U16412 ( .A1(net785255), .A2(n22715), .ZN(n22705) );
  AND2_X1 U16413 ( .A1(net785255), .A2(n22716), .ZN(n22706) );
  AND2_X1 U16414 ( .A1(net785255), .A2(n22710), .ZN(n22707) );
  INV_X1 U16415 ( .A(n26528), .ZN(n22712) );
  INV_X1 U16416 ( .A(n22721), .ZN(n22720) );
  NAND2_X1 U16417 ( .A1(n22708), .A2(n22874), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_23/N3 ) );
  NAND2_X1 U16418 ( .A1(net742649), .A2(n22709), .ZN(n22708) );
  NOR2_X1 U16419 ( .A1(n24582), .A2(n26705), .ZN(n22709) );
  INV_X1 U16420 ( .A(n26382), .ZN(n22711) );
  NAND2_X1 U16421 ( .A1(n22689), .A2(n22711), .ZN(n22710) );
  NAND2_X1 U16422 ( .A1(net716385), .A2(n22712), .ZN(n22713) );
  NAND2_X1 U16423 ( .A1(n22713), .A2(n26527), .ZN(n22714) );
  CLKBUF_X3 U16424 ( .A(net716339), .Z(net796193) );
  CLKBUF_X3 U16425 ( .A(net716339), .Z(net716311) );
  NAND2_X1 U16426 ( .A1(n22690), .A2(n22670), .ZN(n22715) );
  NAND2_X1 U16427 ( .A1(n22691), .A2(n22671), .ZN(n22716) );
  NAND2_X1 U16428 ( .A1(n22717), .A2(n26672), .ZN(
        \core_inst/IF_stage/PROGRAM_COUNTER/DFF_10/N3 ) );
  OR2_X1 U16429 ( .A1(net716387), .A2(n26739), .ZN(n22717) );
  NAND2_X1 U16430 ( .A1(n22718), .A2(n22722), .ZN(n22719) );
  NAND2_X1 U16431 ( .A1(net742576), .A2(n22720), .ZN(n22718) );
  CLKBUF_X3 U16432 ( .A(net716339), .Z(net716313) );
  OAI21_X1 U16433 ( .B1(n22723), .B2(n22724), .A(net717052), .ZN(n22721) );
  NAND4_X1 U16434 ( .A1(n18814), .A2(n22729), .A3(n18815), .A4(n22727), .ZN(
        n22723) );
  AND3_X1 U16435 ( .A1(n18828), .A2(n18827), .A3(n18826), .ZN(n22729) );
  AND2_X1 U16436 ( .A1(n18817), .A2(n18816), .ZN(n22727) );
  NAND4_X1 U16437 ( .A1(n22728), .A2(n18833), .A3(n18825), .A4(n18832), .ZN(
        n22724) );
  AND3_X1 U16438 ( .A1(n18831), .A2(n22725), .A3(n22726), .ZN(n22728) );
  OR2_X1 U16439 ( .A1(n18332), .A2(n818), .ZN(n22725) );
  NAND2_X1 U16440 ( .A1(net767238), .A2(net741400), .ZN(n22726) );
  INV_X1 U16441 ( .A(net767169), .ZN(net767238) );
  BUF_X1 U16442 ( .A(n18326), .Z(net716417) );
  NAND3_X1 U16443 ( .A1(net796255), .A2(net712397), .A3(net712645), .ZN(n22722) );
  AND2_X1 U16444 ( .A1(net713412), .A2(net713413), .ZN(net712397) );
  INV_X1 U16445 ( .A(net717153), .ZN(net712645) );
  NAND2_X1 U16446 ( .A1(net712499), .A2(net712645), .ZN(net795259) );
  NAND3_X1 U16447 ( .A1(net713389), .A2(net713424), .A3(net713425), .ZN(
        net713412) );
  INV_X1 U16448 ( .A(net713414), .ZN(net713413) );
  AND2_X1 U16449 ( .A1(net715884), .A2(net715885), .ZN(net717153) );
  AND2_X1 U16450 ( .A1(net713412), .A2(net713413), .ZN(net717050) );
  AND2_X1 U16451 ( .A1(net716257), .A2(net794712), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_21/N3 ) );
  AND2_X1 U16452 ( .A1(net716257), .A2(n22682), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_31/N3 ) );
  AND2_X1 U16453 ( .A1(net716263), .A2(n22855), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_30/N3 ) );
  AND2_X1 U16454 ( .A1(net716257), .A2(n14195), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_2/N3 ) );
  AND2_X1 U16455 ( .A1(net716253), .A2(n22734), .ZN(n22730) );
  AND2_X1 U16456 ( .A1(net716243), .A2(n22733), .ZN(n22731) );
  NOR2_X1 U16457 ( .A1(net812952), .A2(n23272), .ZN(n23981) );
  NAND2_X1 U16458 ( .A1(net716265), .A2(net741345), .ZN(
        \core_inst/EXMEM_IR/DFF_31/data_reg/n15 ) );
  AND2_X1 U16459 ( .A1(net716257), .A2(n22732), .ZN(
        \core_inst/IDEX_NPC/DFF_0/N3 ) );
  BUF_X2 U16460 ( .A(n15091), .Z(net716385) );
  INV_X1 U16461 ( .A(net765318), .ZN(net826165) );
  OR2_X1 U16462 ( .A1(n26507), .A2(n26506), .ZN(n22733) );
  CLKBUF_X1 U16463 ( .A(net716337), .Z(net796156) );
  OR2_X1 U16464 ( .A1(n26591), .A2(n26590), .ZN(n22734) );
  AND2_X1 U16465 ( .A1(net742612), .A2(n22735), .ZN(
        \core_inst/IDEX_RF_IN1/DFF_7/N3 ) );
  NAND2_X1 U16466 ( .A1(n26677), .A2(n26676), .ZN(n22735) );
  INV_X1 U16467 ( .A(net716385), .ZN(net812958) );
  AND2_X1 U16468 ( .A1(net716263), .A2(n22745), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_8/N3 ) );
  INV_X1 U16469 ( .A(net742612), .ZN(net812952) );
  AND2_X1 U16470 ( .A1(net716263), .A2(n22736), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_14/N3 ) );
  AND2_X1 U16471 ( .A1(net716385), .A2(n22737), .ZN(
        \core_inst/IDEX_RF_IN1/DFF_12/N3 ) );
  NAND2_X1 U16472 ( .A1(n26668), .A2(n26667), .ZN(n22737) );
  INV_X1 U16473 ( .A(net795993), .ZN(net812941) );
  OR2_X2 U16474 ( .A1(net716341), .A2(n23536), .ZN(n24261) );
  OR2_X1 U16475 ( .A1(n24273), .A2(n23611), .ZN(n22738) );
  AND2_X1 U16476 ( .A1(net716263), .A2(n24123), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_23/N3 ) );
  AND2_X1 U16477 ( .A1(net765341), .A2(n22940), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_29/N3 ) );
  OR4_X1 U16478 ( .A1(n23104), .A2(n26567), .A3(net712857), .A4(net712856), 
        .ZN(n22940) );
  BUF_X2 U16479 ( .A(n15091), .Z(net742576) );
  NOR2_X1 U16480 ( .A1(net716353), .A2(n22739), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_31/N3 ) );
  AND2_X1 U16481 ( .A1(net716259), .A2(s_IFID_IR[19]), .ZN(n22740) );
  INV_X1 U16482 ( .A(net712391), .ZN(net812866) );
  BUF_X1 U16483 ( .A(n15091), .Z(net765318) );
  AND3_X2 U16484 ( .A1(net749368), .A2(net731203), .A3(net714705), .ZN(
        net717564) );
  INV_X1 U16486 ( .A(net765318), .ZN(net812284) );
  BUF_X1 U16487 ( .A(net717950), .Z(net795568) );
  INV_X1 U16488 ( .A(net716387), .ZN(net812279) );
  NAND2_X1 U16489 ( .A1(net765318), .A2(net780181), .ZN(n22742) );
  NAND2_X1 U16490 ( .A1(net716387), .A2(net780181), .ZN(net755061) );
  INV_X1 U16491 ( .A(n24284), .ZN(n22745) );
  NAND2_X1 U16497 ( .A1(net716249), .A2(n22681), .ZN(n26350) );
  INV_X1 U16505 ( .A(net712359), .ZN(n22759) );
  NOR2_X1 U16506 ( .A1(net749609), .A2(net720496), .ZN(net742051) );
  NOR2_X1 U16507 ( .A1(net715785), .A2(net715786), .ZN(net749609) );
  NOR2_X1 U16508 ( .A1(net720497), .A2(net715746), .ZN(net720496) );
  NOR2_X1 U16509 ( .A1(net742051), .A2(net717802), .ZN(net715432) );
  NOR2_X1 U16510 ( .A1(net742051), .A2(net742012), .ZN(net717720) );
  NOR2_X1 U16511 ( .A1(net715770), .A2(net89524), .ZN(net715774) );
  NOR2_X1 U16512 ( .A1(net715614), .A2(net720496), .ZN(net715632) );
  AND2_X2 U16513 ( .A1(net742012), .A2(net749609), .ZN(net715445) );
  OR2_X1 U16514 ( .A1(net715747), .A2(net715746), .ZN(net727275) );
  CLKBUF_X1 U16515 ( .A(net742288), .Z(net742282) );
  NAND3_X1 U16516 ( .A1(net715787), .A2(net742288), .A3(net715751), .ZN(
        net715786) );
  INV_X1 U16517 ( .A(net715774), .ZN(net715772) );
  NOR3_X1 U16518 ( .A1(net715774), .A2(net755063), .A3(net715773), .ZN(
        net715787) );
  NAND2_X1 U16519 ( .A1(net715591), .A2(net718092), .ZN(net715785) );
  NAND2_X1 U16520 ( .A1(net742011), .A2(net715661), .ZN(net715751) );
  AOI22_X1 U16521 ( .A1(net750145), .A2(net89524), .B1(net715769), .B2(
        net741339), .ZN(net786871) );
  NAND3_X1 U16522 ( .A1(net804458), .A2(net720724), .A3(net749829), .ZN(
        net715770) );
  NOR2_X1 U16523 ( .A1(net715786), .A2(net715785), .ZN(net715614) );
  AND2_X1 U16524 ( .A1(net715751), .A2(net718092), .ZN(net773963) );
  BUF_X1 U16525 ( .A(net786871), .Z(net717843) );
  NAND2_X1 U16526 ( .A1(net715770), .A2(net715788), .ZN(net715661) );
  AOI22_X1 U16527 ( .A1(net715799), .A2(net89524), .B1(net715769), .B2(
        net741339), .ZN(net715692) );
  NAND2_X1 U16528 ( .A1(net713695), .A2(net715167), .ZN(net714323) );
  INV_X1 U16529 ( .A(net713749), .ZN(net713695) );
  XNOR2_X1 U16530 ( .A(net714961), .B(net716215), .ZN(net715167) );
  NAND2_X1 U16531 ( .A1(net715170), .A2(net715169), .ZN(net714961) );
  INV_X4 U16532 ( .A(net741307), .ZN(net716215) );
  NAND2_X1 U16533 ( .A1(net720607), .A2(net714323), .ZN(net749831) );
  NAND2_X1 U16534 ( .A1(net714323), .A2(net720607), .ZN(net714742) );
  MUX2_X1 U16535 ( .A(net714058), .B(n5582), .S(net741686), .Z(net713749) );
  CLKBUF_X1 U16536 ( .A(net713695), .Z(net755134) );
  NOR3_X1 U16537 ( .A1(n22762), .A2(n22760), .A3(n22761), .ZN(net714058) );
  BUF_X1 U16538 ( .A(net713749), .Z(net718372) );
  OAI22_X1 U16539 ( .A1(net718336), .A2(n17893), .B1(net717719), .B2(n4331), 
        .ZN(n22762) );
  INV_X1 U16540 ( .A(net715445), .ZN(net718336) );
  INV_X1 U16541 ( .A(net715432), .ZN(net717719) );
  NOR2_X1 U16542 ( .A1(net717594), .A2(n5609), .ZN(n22760) );
  INV_X1 U16543 ( .A(net742284), .ZN(net717594) );
  AND2_X1 U16544 ( .A1(net750018), .A2(\core_inst/MEMWB_ALUOUT/DFF_8/N3 ), 
        .ZN(n22761) );
  CLKBUF_X1 U16545 ( .A(net750135), .Z(net750018) );
  MUX2_X1 U16546 ( .A(n5582), .B(net714058), .S(net787526), .Z(net786844) );
  CLKBUF_X1 U16547 ( .A(net714058), .Z(net742042) );
  NAND2_X1 U16548 ( .A1(net727275), .A2(net715748), .ZN(net717802) );
  BUF_X1 U16549 ( .A(net715432), .Z(net742265) );
  INV_X1 U16550 ( .A(net715432), .ZN(net717718) );
  OAI22_X1 U16551 ( .A1(net718336), .A2(net740717), .B1(net715419), .B2(n1696), 
        .ZN(net768639) );
  OAI22_X1 U16552 ( .A1(n4347), .A2(net718336), .B1(net742413), .B2(n1752), 
        .ZN(net715576) );
  OAI22_X1 U16553 ( .A1(n1736), .A2(net718432), .B1(net740721), .B2(net718336), 
        .ZN(net715418) );
  AOI22_X1 U16554 ( .A1(net741609), .A2(net741580), .B1(net741527), .B2(
        net741293), .ZN(net715847) );
  OAI22_X1 U16555 ( .A1(n1726), .A2(net749972), .B1(net714943), .B2(n17893), 
        .ZN(net715171) );
  NOR2_X1 U16556 ( .A1(net762680), .A2(n4331), .ZN(net715172) );
  AND2_X2 U16557 ( .A1(net717802), .A2(net715615), .ZN(net750135) );
  BUF_X2 U16558 ( .A(net717802), .Z(net749369) );
  OAI21_X1 U16559 ( .B1(net773962), .B2(net773961), .A(net773963), .ZN(
        net715748) );
  XNOR2_X1 U16560 ( .A(net714961), .B(net716231), .ZN(net750182) );
  OAI22_X1 U16561 ( .A1(n5589), .A2(net717594), .B1(net717718), .B2(n4352), 
        .ZN(net715598) );
  OAI22_X1 U16562 ( .A1(net717594), .A2(net740634), .B1(n4409), .B2(net717719), 
        .ZN(net715551) );
  OAI22_X1 U16563 ( .A1(net717594), .A2(net740632), .B1(net717718), .B2(n4388), 
        .ZN(net747437) );
  AOI22_X1 U16564 ( .A1(net750018), .A2(\core_inst/MEMWB_ALUOUT/DFF_24/N3 ), 
        .B1(net750111), .B2(n640), .ZN(net715536) );
  AND2_X1 U16565 ( .A1(net715748), .A2(net727275), .ZN(net737672) );
  NAND2_X1 U16566 ( .A1(net727275), .A2(net715748), .ZN(net742012) );
  OAI211_X1 U16567 ( .C1(n22769), .C2(n22766), .A(n22770), .B(n22767), .ZN(
        net738752) );
  OR2_X1 U16568 ( .A1(net717607), .A2(net760174), .ZN(n22769) );
  AND2_X1 U16569 ( .A1(net713921), .A2(net717564), .ZN(net717607) );
  AND2_X1 U16570 ( .A1(net755215), .A2(net713905), .ZN(net760174) );
  NAND2_X1 U16571 ( .A1(net727668), .A2(net749633), .ZN(n22766) );
  AND3_X1 U16572 ( .A1(n22772), .A2(n22773), .A3(n22774), .ZN(n22770) );
  NAND3_X1 U16573 ( .A1(net780581), .A2(net749830), .A3(n22771), .ZN(n22772)
         );
  NOR2_X1 U16574 ( .A1(net732820), .A2(net732819), .ZN(net780581) );
  AND3_X1 U16575 ( .A1(net713833), .A2(net714705), .A3(net731203), .ZN(
        net749830) );
  AND2_X1 U16576 ( .A1(net735179), .A2(net760174), .ZN(n22771) );
  NOR2_X1 U16577 ( .A1(net713924), .A2(net713154), .ZN(n22773) );
  INV_X1 U16578 ( .A(net714544), .ZN(net713924) );
  INV_X2 U16579 ( .A(net712459), .ZN(net713154) );
  NAND2_X1 U16580 ( .A1(net712880), .A2(n22768), .ZN(n22774) );
  NAND2_X1 U16581 ( .A1(net713966), .A2(net714934), .ZN(net712880) );
  INV_X1 U16582 ( .A(net760174), .ZN(n22768) );
  NAND2_X1 U16583 ( .A1(n22766), .A2(n22771), .ZN(n22767) );
  NAND2_X1 U16584 ( .A1(net738752), .A2(net738751), .ZN(net736102) );
  NOR2_X1 U16585 ( .A1(net732819), .A2(net732820), .ZN(net713921) );
  NOR2_X1 U16586 ( .A1(n22764), .A2(n22763), .ZN(net732819) );
  NAND2_X1 U16587 ( .A1(net714702), .A2(net736222), .ZN(net732820) );
  OR2_X1 U16588 ( .A1(net725613), .A2(net717607), .ZN(net713806) );
  INV_X1 U16589 ( .A(net717607), .ZN(net749400) );
  OAI21_X1 U16590 ( .B1(net714703), .B2(net742308), .A(net740525), .ZN(n22764)
         );
  NAND2_X1 U16591 ( .A1(net714856), .A2(net714136), .ZN(net714703) );
  AND2_X2 U16592 ( .A1(net714742), .A2(net714749), .ZN(net742308) );
  NAND2_X1 U16593 ( .A1(net762630), .A2(net714833), .ZN(net740525) );
  NOR3_X1 U16594 ( .A1(n22765), .A2(net742308), .A3(net767320), .ZN(n22763) );
  OAI21_X1 U16595 ( .B1(net742146), .B2(net755139), .A(net714860), .ZN(n22765)
         );
  OR2_X2 U16596 ( .A1(net755210), .A2(net713754), .ZN(net742146) );
  XNOR2_X1 U16597 ( .A(net749698), .B(net716231), .ZN(net755139) );
  INV_X1 U16598 ( .A(net714861), .ZN(net714860) );
  INV_X1 U16599 ( .A(net714975), .ZN(net767320) );
  OR2_X1 U16600 ( .A1(net732820), .A2(net732819), .ZN(net749945) );
  NAND2_X1 U16601 ( .A1(net749831), .A2(net714749), .ZN(net762630) );
  NAND2_X1 U16602 ( .A1(net713709), .A2(net753295), .ZN(net714749) );
  NAND2_X1 U16603 ( .A1(net714328), .A2(net714749), .ZN(net714833) );
  CLKBUF_X1 U16604 ( .A(net740525), .Z(net755097) );
  NAND2_X1 U16605 ( .A1(net755642), .A2(net783365), .ZN(net720607) );
  NAND2_X1 U16606 ( .A1(net749831), .A2(net714749), .ZN(net714128) );
  NOR2_X1 U16607 ( .A1(net714539), .A2(net760174), .ZN(net714545) );
  INV_X1 U16608 ( .A(net717564), .ZN(net714113) );
  AND2_X1 U16609 ( .A1(net780581), .A2(net717564), .ZN(net765361) );
  OR2_X1 U16610 ( .A1(net731060), .A2(net717564), .ZN(net713943) );
  NAND3_X1 U16611 ( .A1(net758890), .A2(net714703), .A3(net758891), .ZN(
        net714702) );
  NAND2_X1 U16612 ( .A1(net714703), .A2(net742275), .ZN(net714157) );
  NOR2_X1 U16613 ( .A1(net755086), .A2(net742308), .ZN(net778368) );
  INV_X1 U16614 ( .A(net742308), .ZN(net742286) );
  NOR3_X1 U16615 ( .A1(net746029), .A2(net714833), .A3(net714747), .ZN(
        net714285) );
  NOR2_X1 U16616 ( .A1(net714833), .A2(net714855), .ZN(net758891) );
  AND2_X1 U16617 ( .A1(net714128), .A2(net714833), .ZN(net714551) );
  NAND2_X1 U16618 ( .A1(net717547), .A2(net749428), .ZN(net727668) );
  BUF_X1 U16619 ( .A(net718400), .Z(net749633) );
  XOR2_X1 U16620 ( .A(net713934), .B(net716215), .Z(net755215) );
  INV_X2 U16621 ( .A(net713570), .ZN(net713905) );
  NAND3_X1 U16622 ( .A1(net766153), .A2(net733611), .A3(net739130), .ZN(
        net749368) );
  AND2_X1 U16623 ( .A1(net714709), .A2(net714599), .ZN(net731203) );
  OAI21_X1 U16624 ( .B1(net714706), .B2(net714610), .A(net730300), .ZN(
        net714705) );
  NAND3_X1 U16625 ( .A1(net728823), .A2(net769908), .A3(net728824), .ZN(
        net736222) );
  OAI21_X1 U16626 ( .B1(net780578), .B2(net714858), .A(net749841), .ZN(
        net714856) );
  NAND2_X1 U16627 ( .A1(net749841), .A2(net715032), .ZN(net714136) );
  NAND2_X1 U16628 ( .A1(net718372), .A2(net750182), .ZN(net714328) );
  XNOR2_X1 U16629 ( .A(net713710), .B(net716223), .ZN(net753295) );
  INV_X1 U16630 ( .A(net713709), .ZN(net755642) );
  XNOR2_X1 U16631 ( .A(net713710), .B(net716215), .ZN(net783365) );
  NAND2_X1 U16632 ( .A1(net727668), .A2(net749945), .ZN(net714104) );
  NAND2_X1 U16633 ( .A1(net749476), .A2(net749633), .ZN(net725613) );
  NOR2_X1 U16634 ( .A1(net755215), .A2(net713154), .ZN(net738766) );
  NAND2_X1 U16635 ( .A1(net755215), .A2(net713905), .ZN(net713923) );
  AND2_X1 U16636 ( .A1(net738443), .A2(net749368), .ZN(net749507) );
  OAI21_X1 U16637 ( .B1(net714754), .B2(net714157), .A(net714702), .ZN(
        net714770) );
  INV_X1 U16638 ( .A(net714136), .ZN(net758644) );
  AND2_X1 U16639 ( .A1(net804677), .A2(net714136), .ZN(net746029) );
  CLKBUF_X1 U16640 ( .A(net714742), .Z(net804675) );
  AND2_X1 U16641 ( .A1(net714328), .A2(net714749), .ZN(net742275) );
  CLKBUF_X1 U16642 ( .A(net783365), .Z(net786821) );
  AOI21_X1 U16643 ( .B1(net717091), .B2(net780200), .A(net780201), .ZN(
        net712359) );
  INV_X1 U16644 ( .A(net716337), .ZN(net716243) );
  INV_X1 U16645 ( .A(net712487), .ZN(net712486) );
  NOR2_X1 U16646 ( .A1(net712976), .A2(net760170), .ZN(net713492) );
  OAI21_X1 U16647 ( .B1(net724352), .B2(net724353), .A(net724354), .ZN(
        net712966) );
  OAI211_X1 U16648 ( .C1(net713495), .C2(net712975), .A(net713496), .B(
        net712971), .ZN(net713493) );
  INV_X1 U16649 ( .A(net712965), .ZN(net713494) );
  NOR2_X1 U16650 ( .A1(n22777), .A2(net713758), .ZN(net713757) );
  OAI21_X1 U16651 ( .B1(net712473), .B2(net713154), .A(net712472), .ZN(n22777)
         );
  AOI22_X1 U16652 ( .A1(net713803), .A2(net713804), .B1(net713806), .B2(
        net713805), .ZN(net712473) );
  AOI211_X1 U16653 ( .C1(net713760), .C2(net713761), .A(net713762), .B(
        net713763), .ZN(net712472) );
  NAND2_X1 U16654 ( .A1(net734492), .A2(net726730), .ZN(net726729) );
  XNOR2_X1 U16655 ( .A(net735735), .B(net713995), .ZN(net734492) );
  INV_X1 U16656 ( .A(net712844), .ZN(net726730) );
  NOR2_X1 U16657 ( .A1(net713849), .A2(net713850), .ZN(net713074) );
  NAND3_X1 U16658 ( .A1(net713858), .A2(net713859), .A3(net713860), .ZN(
        net713849) );
  AOI21_X1 U16659 ( .B1(net712462), .B2(net712469), .A(net729186), .ZN(
        net713850) );
  NOR3_X1 U16660 ( .A1(n22778), .A2(net736102), .A3(n22779), .ZN(net713756) );
  NOR2_X1 U16661 ( .A1(n22799), .A2(n22782), .ZN(n22778) );
  AND2_X1 U16662 ( .A1(n22780), .A2(n22781), .ZN(n22799) );
  NOR2_X1 U16663 ( .A1(n22789), .A2(n22790), .ZN(n22780) );
  INV_X1 U16664 ( .A(n22786), .ZN(n22789) );
  OAI21_X1 U16665 ( .B1(net713964), .B2(net755060), .A(net755714), .ZN(n22786)
         );
  NAND2_X1 U16666 ( .A1(n22791), .A2(net713943), .ZN(n22790) );
  INV_X1 U16667 ( .A(n22787), .ZN(n22791) );
  MUX2_X1 U16668 ( .A(net713949), .B(net713951), .S(net713950), .Z(n22787) );
  NAND2_X1 U16669 ( .A1(net713152), .A2(net749936), .ZN(net713949) );
  NAND2_X1 U16670 ( .A1(net713148), .A2(net715351), .ZN(net713951) );
  XNOR2_X1 U16671 ( .A(net713967), .B(net716221), .ZN(net713950) );
  NAND3_X1 U16672 ( .A1(net713952), .A2(net734385), .A3(net713168), .ZN(n22781) );
  OAI21_X1 U16673 ( .B1(n22783), .B2(n22781), .A(n22784), .ZN(n22782) );
  INV_X1 U16674 ( .A(n22788), .ZN(n22783) );
  OAI22_X1 U16675 ( .A1(net713949), .A2(net713829), .B1(net713951), .B2(
        net713950), .ZN(n22788) );
  OAI21_X1 U16676 ( .B1(net713154), .B2(n22788), .A(n22785), .ZN(n22784) );
  NAND3_X1 U16677 ( .A1(net713943), .A2(net717091), .A3(n22786), .ZN(n22785)
         );
  OAI21_X1 U16678 ( .B1(n22776), .B2(net712844), .A(n22775), .ZN(n22779) );
  INV_X1 U16679 ( .A(net713909), .ZN(n22776) );
  NAND2_X1 U16680 ( .A1(net742508), .A2(net713993), .ZN(net713909) );
  OAI22_X1 U16681 ( .A1(net713909), .A2(net717091), .B1(net742507), .B2(
        net713910), .ZN(net712844) );
  INV_X1 U16682 ( .A(net746686), .ZN(n22775) );
  OAI211_X1 U16683 ( .C1(net713857), .C2(net729186), .A(net746687), .B(
        net746688), .ZN(net746686) );
  NOR3_X1 U16684 ( .A1(net712447), .A2(net712840), .A3(net712841), .ZN(
        net713755) );
  AND2_X1 U16685 ( .A1(net749239), .A2(net712459), .ZN(net712447) );
  NOR2_X1 U16686 ( .A1(net734492), .A2(net713992), .ZN(net712840) );
  NAND2_X1 U16687 ( .A1(net713909), .A2(net717091), .ZN(net713992) );
  NAND4_X1 U16688 ( .A1(net713973), .A2(net713974), .A3(net713975), .A4(
        net713976), .ZN(net712841) );
  NAND2_X1 U16689 ( .A1(n22792), .A2(n22793), .ZN(net738751) );
  OAI21_X1 U16690 ( .B1(net765361), .B2(net725613), .A(n22798), .ZN(n22792) );
  NOR2_X1 U16691 ( .A1(net712880), .A2(n22795), .ZN(n22798) );
  NAND2_X1 U16692 ( .A1(net713767), .A2(net713930), .ZN(n22795) );
  INV_X1 U16693 ( .A(n22794), .ZN(n22793) );
  OAI22_X1 U16694 ( .A1(n22795), .A2(net738766), .B1(net746701), .B2(n22796), 
        .ZN(n22794) );
  INV_X1 U16695 ( .A(net713905), .ZN(net746701) );
  OAI21_X1 U16696 ( .B1(net762674), .B2(net713728), .A(n22797), .ZN(n22796) );
  AND3_X1 U16697 ( .A1(net724630), .A2(net724632), .A3(net724631), .ZN(
        net762674) );
  NAND2_X1 U16698 ( .A1(net762674), .A2(net713736), .ZN(n22797) );
  INV_X1 U16699 ( .A(net713770), .ZN(net713736) );
  CLKBUF_X1 U16700 ( .A(net736102), .Z(net749607) );
  NOR2_X1 U16701 ( .A1(net716313), .A2(net712359), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_14/N3 ) );
  OAI21_X1 U16702 ( .B1(net712377), .B2(net716267), .A(net712737), .ZN(
        net522736) );
  AND2_X1 U16703 ( .A1(net716243), .A2(net712486), .ZN(net767257) );
  INV_X1 U16704 ( .A(net712494), .ZN(net780200) );
  INV_X1 U16705 ( .A(net712493), .ZN(net780201) );
  CLKBUF_X1 U16706 ( .A(net716341), .Z(net796133) );
  OAI21_X1 U16707 ( .B1(net712488), .B2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [14]), .A(net712490), .ZN(net712487) );
  CLKBUF_X1 U16708 ( .A(net713492), .Z(net780542) );
  AOI21_X1 U16709 ( .B1(net712966), .B2(net712967), .A(net712968), .ZN(
        net712964) );
  AOI22_X1 U16710 ( .A1(net780542), .A2(net712966), .B1(net785249), .B2(
        net713494), .ZN(net755094) );
  CLKBUF_X1 U16711 ( .A(net713493), .Z(net785249) );
  NOR2_X1 U16712 ( .A1(net712447), .A2(net796127), .ZN(net712376) );
  AOI211_X1 U16713 ( .C1(net726730), .C2(net780215), .A(net712841), .B(
        net795962), .ZN(net712365) );
  CLKBUF_X1 U16714 ( .A(n26112), .Z(n22800) );
  AOI21_X1 U16715 ( .B1(n23931), .B2(net714858), .A(n24040), .ZN(net804677) );
  NOR2_X2 U16716 ( .A1(n23576), .A2(n25576), .ZN(net714858) );
  AND2_X1 U16717 ( .A1(net765341), .A2(n22802), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_23/N3 ) );
  AOI21_X1 U16718 ( .B1(n22804), .B2(n22805), .A(net796143), .ZN(n22803) );
  OR2_X1 U16719 ( .A1(n24008), .A2(n23067), .ZN(n22804) );
  NAND2_X1 U16720 ( .A1(net717050), .A2(n26662), .ZN(n22805) );
  AOI21_X1 U16721 ( .B1(n22807), .B2(n22808), .A(net796232), .ZN(n22806) );
  OR2_X1 U16722 ( .A1(n26637), .A2(n26358), .ZN(n22807) );
  NAND2_X1 U16723 ( .A1(net717048), .A2(n26436), .ZN(n22808) );
  NOR2_X1 U16724 ( .A1(net812941), .A2(n22809), .ZN(
        \core_inst/IFID_IR/DFF_21/N3 ) );
  INV_X32 U16725 ( .A(\core_inst/s_IF_OUT_IR_OUT [21]), .ZN(n22809) );
  INV_X1 U16726 ( .A(net716265), .ZN(net804641) );
  INV_X1 U16727 ( .A(n26569), .ZN(n22810) );
  NOR2_X1 U16728 ( .A1(net765319), .A2(n22811), .ZN(
        \core_inst/EXMEM_RF_ADDR_DEST/DFF_1/N3 ) );
  INV_X1 U16729 ( .A(n24156), .ZN(n22812) );
  AOI22_X1 U16730 ( .A1(n22850), .A2(n24362), .B1(n24363), .B2(n24364), .ZN(
        n22813) );
  CLKBUF_X1 U16731 ( .A(n26231), .Z(n23381) );
  AND2_X1 U16732 ( .A1(net760161), .A2(n22814), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_17/N3 ) );
  AND2_X1 U16733 ( .A1(net716259), .A2(n23513), .ZN(n22815) );
  AND2_X1 U16734 ( .A1(net716385), .A2(n25336), .ZN(n26742) );
  NAND2_X1 U16735 ( .A1(net765341), .A2(n22816), .ZN(n23946) );
  CLKBUF_X3 U16736 ( .A(net716339), .Z(net716333) );
  INV_X1 U16737 ( .A(net742576), .ZN(net804592) );
  CLKBUF_X1 U16738 ( .A(net718092), .Z(net750053) );
  CLKBUF_X1 U16739 ( .A(n24320), .Z(n24193) );
  INV_X1 U16740 ( .A(n26703), .ZN(n22832) );
  OAI22_X1 U16741 ( .A1(net715058), .A2(n25321), .B1(net738474), .B2(n1628), 
        .ZN(n23723) );
  NAND2_X1 U16742 ( .A1(n22820), .A2(n22817), .ZN(net804458) );
  NOR2_X1 U16743 ( .A1(net741237), .A2(net741262), .ZN(n22817) );
  NAND2_X1 U16744 ( .A1(net720730), .A2(net741345), .ZN(net720724) );
  NAND2_X1 U16745 ( .A1(net720729), .A2(net720728), .ZN(net749829) );
  NAND2_X1 U16746 ( .A1(n14130), .A2(n14382), .ZN(net720729) );
  NOR2_X1 U16747 ( .A1(n15079), .A2(n14073), .ZN(net720728) );
  XNOR2_X1 U16748 ( .A(net718078), .B(net718077), .ZN(n22820) );
  NAND3_X1 U16749 ( .A1(net804458), .A2(net720725), .A3(net720724), .ZN(
        net742011) );
  NOR2_X1 U16750 ( .A1(net716313), .A2(net741262), .ZN(
        \core_inst/EXMEM_IR/DFF_27/N3 ) );
  NAND3_X1 U16751 ( .A1(net741262), .A2(n14073), .A3(net749566), .ZN(n22818)
         );
  NAND3_X1 U16752 ( .A1(n15079), .A2(net741576), .A3(net741237), .ZN(n22819)
         );
  BUF_X1 U16753 ( .A(n14130), .Z(net749566) );
  OR2_X1 U16754 ( .A1(net718078), .A2(net718077), .ZN(net720730) );
  INV_X1 U16755 ( .A(n14389), .ZN(net715790) );
  AND2_X1 U16756 ( .A1(net742648), .A2(n14389), .ZN(
        \core_inst/EXMEM_IR/DFF_30/N3 ) );
  NAND4_X1 U16757 ( .A1(n22818), .A2(net715790), .A3(n22819), .A4(net741345), 
        .ZN(net715788) );
  NAND2_X1 U16758 ( .A1(net720729), .A2(net720728), .ZN(net720725) );
  OAI211_X1 U16759 ( .C1(net714743), .C2(net804675), .A(net714744), .B(
        net718140), .ZN(net714164) );
  OAI211_X1 U16760 ( .C1(net812773), .C2(n13165), .A(n22821), .B(net755061), 
        .ZN(\core_inst/IDEX_RF_ADDR_DEST/DFF_1/N3 ) );
  NAND2_X1 U16761 ( .A1(n22822), .A2(s_IFID_IR[17]), .ZN(n22821) );
  NOR2_X1 U16762 ( .A1(net713485), .A2(net795568), .ZN(n22822) );
  NOR3_X1 U16763 ( .A1(n18137), .A2(net710357), .A3(n18130), .ZN(net713485) );
  NAND2_X1 U16764 ( .A1(n22822), .A2(s_IFID_IR[19]), .ZN(net713484) );
  NAND2_X1 U16765 ( .A1(n22822), .A2(s_IFID_IR[20]), .ZN(net713480) );
  OAI211_X1 U16766 ( .C1(net812773), .C2(n6562), .A(net713484), .B(net755061), 
        .ZN(\core_inst/IDEX_RF_ADDR_DEST/DFF_3/N3 ) );
  NOR2_X1 U16767 ( .A1(net796200), .A2(n13165), .ZN(net712313) );
  INV_X1 U16768 ( .A(net713485), .ZN(net718074) );
  NAND2_X1 U16769 ( .A1(net713389), .A2(net518455), .ZN(n18136) );
  BUF_X1 U16770 ( .A(n15091), .Z(net795993) );
  AND2_X1 U16771 ( .A1(net718074), .A2(n18136), .ZN(net780181) );
  NAND3_X1 U16772 ( .A1(n20115), .A2(net709330), .A3(n18158), .ZN(n18137) );
  INV_X1 U16773 ( .A(net518455), .ZN(net710357) );
  INV_X1 U16774 ( .A(n18135), .ZN(n18130) );
  NOR3_X1 U16775 ( .A1(n18137), .A2(n18130), .A3(net741279), .ZN(net710387) );
  AOI211_X1 U16776 ( .C1(net710357), .C2(s_IFID_IR[30]), .A(n18143), .B(n18196), .ZN(n20115) );
  NOR4_X1 U16777 ( .A1(n18130), .A2(net712961), .A3(net720303), .A4(net720304), 
        .ZN(net720302) );
  NAND2_X1 U16778 ( .A1(net742368), .A2(n22679), .ZN(n25550) );
  CLKBUF_X1 U16779 ( .A(net716337), .Z(net796271) );
  MUX2_X1 U16780 ( .A(\core_inst/EXMEM_NPC/DFF_14/N3 ), .B(n26091), .S(
        net716237), .Z(n24548) );
  INV_X1 U16781 ( .A(net713733), .ZN(net796258) );
  AND3_X2 U16782 ( .A1(n23751), .A2(n23750), .A3(n23749), .ZN(n24381) );
  AND2_X1 U16783 ( .A1(net760161), .A2(n22823), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_10/N3 ) );
  AND2_X1 U16784 ( .A1(net760161), .A2(\core_inst/s_IF_OUT_IR_OUT [29]), .ZN(
        \core_inst/IFID_IR/DFF_29/N3 ) );
  AND2_X1 U16785 ( .A1(net785255), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/CLA_PG_NET/N1 ), .ZN(
        n22824) );
  AOI21_X1 U16786 ( .B1(n22826), .B2(n22827), .A(net796133), .ZN(n22825) );
  OR2_X1 U16787 ( .A1(n26637), .A2(n26456), .ZN(n22826) );
  NAND2_X1 U16788 ( .A1(n25665), .A2(n26652), .ZN(n22827) );
  AND2_X1 U16789 ( .A1(net716257), .A2(net754762), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_24/N3 ) );
  NOR2_X1 U16790 ( .A1(n24527), .A2(net716311), .ZN(n22828) );
  AND2_X1 U16791 ( .A1(n23538), .A2(n23537), .ZN(n22829) );
  CLKBUF_X1 U16792 ( .A(n26253), .Z(n22830) );
  AOI21_X1 U16793 ( .B1(n23658), .B2(n26213), .A(n26214), .ZN(n26253) );
  XNOR2_X1 U16794 ( .A(n26001), .B(net716223), .ZN(n25872) );
  CLKBUF_X3 U16795 ( .A(net712470), .Z(net796212) );
  AOI21_X1 U16796 ( .B1(n22832), .B2(n22833), .A(net796156), .ZN(n22831) );
  NAND2_X1 U16797 ( .A1(net717050), .A2(n26702), .ZN(n22833) );
  OR2_X1 U16798 ( .A1(net715365), .A2(n24267), .ZN(n26063) );
  CLKBUF_X1 U16799 ( .A(n25425), .Z(n22834) );
  CLKBUF_X1 U16800 ( .A(net716339), .Z(net796200) );
  OAI21_X1 U16801 ( .B1(n23949), .B2(net714610), .A(net730300), .ZN(n22835) );
  CLKBUF_X1 U16802 ( .A(n25780), .Z(n22836) );
  BUF_X1 U16803 ( .A(net731344), .Z(net750024) );
  NOR2_X1 U16804 ( .A1(n23687), .A2(n24549), .ZN(n22837) );
  CLKBUF_X1 U16805 ( .A(n25450), .Z(n24337) );
  AND2_X2 U16806 ( .A1(n24380), .A2(n24381), .ZN(net749843) );
  CLKBUF_X1 U16807 ( .A(net737937), .Z(net796126) );
  NOR2_X2 U16808 ( .A1(n26671), .A2(n5576), .ZN(n26572) );
  NOR2_X2 U16809 ( .A1(n26578), .A2(n6511), .ZN(net712922) );
  NOR2_X2 U16810 ( .A1(n26573), .A2(n11848), .ZN(net712488) );
  NOR2_X2 U16811 ( .A1(net712490), .A2(n6516), .ZN(n26579) );
  AND3_X1 U16812 ( .A1(net742257), .A2(net765400), .A3(net750053), .ZN(
        net796159) );
  AND2_X1 U16813 ( .A1(n22738), .A2(net749289), .ZN(n22838) );
  AOI221_X1 U16814 ( .B1(net749707), .B2(net712872), .C1(n22838), .C2(
        net712872), .A(n24089), .ZN(n23096) );
  NOR2_X1 U16815 ( .A1(net716311), .A2(n22839), .ZN(
        \core_inst/IFID_IR/DFF_23/N3 ) );
  INV_X32 U16816 ( .A(\core_inst/s_IF_OUT_IR_OUT [23]), .ZN(n22839) );
  AND2_X1 U16817 ( .A1(net716255), .A2(net712793), .ZN(n22840) );
  AND2_X1 U16818 ( .A1(net716253), .A2(n22866), .ZN(n22841) );
  AND2_X1 U16819 ( .A1(net760161), .A2(n14190), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_0/N3 ) );
  AND2_X1 U16820 ( .A1(net760161), .A2(s_IFID_IR[26]), .ZN(
        \core_inst/IDEX_IR/DFF_26/N3 ) );
  NOR2_X1 U16821 ( .A1(net765727), .A2(n22842), .ZN(
        \core_inst/IFID_IR/DFF_14/N3 ) );
  INV_X32 U16822 ( .A(\core_inst/s_IF_OUT_IR_OUT [14]), .ZN(n22842) );
  AND2_X1 U16823 ( .A1(net760161), .A2(n23465), .ZN(n22843) );
  INV_X1 U16824 ( .A(net716387), .ZN(net796137) );
  INV_X1 U16825 ( .A(net795993), .ZN(net796136) );
  OR2_X1 U16826 ( .A1(n23963), .A2(n23965), .ZN(n23961) );
  AND2_X1 U16827 ( .A1(n24332), .A2(n23896), .ZN(n22844) );
  BUF_X1 U16828 ( .A(n26131), .Z(n23896) );
  CLKBUF_X1 U16829 ( .A(net746686), .Z(net796127) );
  INV_X1 U16830 ( .A(net717876), .ZN(net796122) );
  BUF_X1 U16831 ( .A(net715632), .Z(net717876) );
  INV_X1 U16832 ( .A(net716387), .ZN(net796114) );
  CLKBUF_X3 U16833 ( .A(net712470), .Z(net717074) );
  MUX2_X2 U16834 ( .A(n829), .B(n26105), .S(net787528), .Z(n26209) );
  XNOR2_X1 U16835 ( .A(n25832), .B(net716215), .ZN(n22845) );
  INV_X1 U16836 ( .A(net714248), .ZN(net796014) );
  OAI211_X1 U16837 ( .C1(n23960), .C2(n23951), .A(n23961), .B(n23962), .ZN(
        n23959) );
  OAI22_X1 U16838 ( .A1(n23017), .A2(net729186), .B1(n23021), .B2(net714382), 
        .ZN(net714415) );
  OAI22_X1 U16839 ( .A1(net749443), .A2(n4391), .B1(net718432), .B2(n1722), 
        .ZN(n25441) );
  NOR2_X1 U16840 ( .A1(net734493), .A2(net713992), .ZN(net795962) );
  OR2_X1 U16842 ( .A1(net716341), .A2(n23544), .ZN(n26708) );
  OR2_X2 U16843 ( .A1(n26239), .A2(n26234), .ZN(n22847) );
  INV_X4 U16844 ( .A(n22847), .ZN(n26242) );
  NAND2_X1 U16846 ( .A1(net716255), .A2(n22680), .ZN(n24077) );
  AND3_X1 U16847 ( .A1(n23605), .A2(n23606), .A3(n23607), .ZN(n22850) );
  CLKBUF_X1 U16848 ( .A(net712976), .Z(net795273) );
  NOR2_X1 U16849 ( .A1(n23768), .A2(n23769), .ZN(n22851) );
  NOR2_X1 U16850 ( .A1(n23768), .A2(n23769), .ZN(n24396) );
  NAND2_X1 U16851 ( .A1(net796255), .A2(n22683), .ZN(n23216) );
  MUX2_X2 U16852 ( .A(\core_inst/EXMEM_NPC/DFF_26/N3 ), .B(n26084), .S(
        net716237), .Z(net713570) );
  AOI21_X1 U16853 ( .B1(n22853), .B2(net795259), .A(net796143), .ZN(n22852) );
  OR2_X1 U16854 ( .A1(n26637), .A2(n26455), .ZN(n22853) );
  INV_X1 U16855 ( .A(net716341), .ZN(net785255) );
  INV_X1 U16857 ( .A(n26727), .ZN(n22856) );
  INV_X1 U16859 ( .A(net712376), .ZN(net794712) );
  OAI22_X1 U16860 ( .A1(net735736), .A2(net735737), .B1(net735738), .B2(
        net748854), .ZN(net735735) );
  NAND2_X1 U16861 ( .A1(n22861), .A2(n22860), .ZN(net735736) );
  NOR2_X1 U16862 ( .A1(n22859), .A2(net720372), .ZN(n22861) );
  NOR2_X1 U16863 ( .A1(n22858), .A2(net714285), .ZN(n22859) );
  NAND3_X1 U16864 ( .A1(net717591), .A2(net767213), .A3(net718140), .ZN(
        net720372) );
  NAND2_X1 U16865 ( .A1(n22862), .A2(n22863), .ZN(n22860) );
  NAND2_X1 U16866 ( .A1(net714006), .A2(net714007), .ZN(n22862) );
  INV_X1 U16867 ( .A(net742309), .ZN(n22863) );
  NOR2_X1 U16868 ( .A1(net714008), .A2(net725077), .ZN(net735737) );
  NAND2_X1 U16869 ( .A1(net714281), .A2(net755735), .ZN(net714008) );
  INV_X1 U16870 ( .A(net713468), .ZN(net725077) );
  NOR3_X1 U16871 ( .A1(n22865), .A2(n22864), .A3(net714002), .ZN(net735738) );
  AOI21_X1 U16872 ( .B1(net714947), .B2(net728158), .A(net714724), .ZN(n22865)
         );
  NAND2_X1 U16873 ( .A1(net714612), .A2(net714611), .ZN(net714947) );
  INV_X1 U16874 ( .A(net714610), .ZN(net728158) );
  INV_X1 U16875 ( .A(net755733), .ZN(net714724) );
  INV_X1 U16876 ( .A(n22863), .ZN(n22864) );
  NAND2_X1 U16877 ( .A1(net749338), .A2(net749905), .ZN(net714002) );
  AND2_X1 U16878 ( .A1(n22862), .A2(n22863), .ZN(net748854) );
  INV_X1 U16879 ( .A(net715146), .ZN(net713995) );
  CLKBUF_X1 U16880 ( .A(net734492), .Z(net734493) );
  OAI21_X1 U16881 ( .B1(net714128), .B2(net714747), .A(net714748), .ZN(n22858)
         );
  INV_X1 U16882 ( .A(n22859), .ZN(net714907) );
  NOR2_X1 U16883 ( .A1(n22859), .A2(net720372), .ZN(net742423) );
  NAND2_X1 U16884 ( .A1(net714119), .A2(net750235), .ZN(net714747) );
  AOI21_X1 U16885 ( .B1(net714439), .B2(net750235), .A(net714842), .ZN(
        net714748) );
  INV_X1 U16886 ( .A(n22858), .ZN(net713468) );
  NOR2_X1 U16887 ( .A1(net714287), .A2(n22858), .ZN(net714950) );
  NOR2_X1 U16888 ( .A1(net713995), .A2(net742507), .ZN(net714586) );
  NOR2_X1 U16889 ( .A1(net713995), .A2(net742508), .ZN(net749542) );
  NAND2_X1 U16890 ( .A1(net720372), .A2(net766652), .ZN(net720121) );
  INV_X1 U16891 ( .A(net720372), .ZN(net734346) );
  CLKBUF_X1 U16892 ( .A(net714285), .Z(net741987) );
  OAI21_X1 U16893 ( .B1(net714746), .B2(net714747), .A(net714748), .ZN(
        net714744) );
  INV_X1 U16894 ( .A(net714748), .ZN(net714743) );
  XNOR2_X1 U16895 ( .A(net713561), .B(net716215), .ZN(net715146) );
  NOR2_X1 U16896 ( .A1(net714751), .A2(net718103), .ZN(net717591) );
  CLKBUF_X2 U16897 ( .A(net755733), .Z(net767213) );
  AND2_X2 U16898 ( .A1(net715050), .A2(net749798), .ZN(net718140) );
  NAND2_X1 U16899 ( .A1(net714440), .A2(net742325), .ZN(net714119) );
  NAND2_X1 U16900 ( .A1(net714123), .A2(net765546), .ZN(net750235) );
  NOR2_X1 U16901 ( .A1(net714440), .A2(net742325), .ZN(net714439) );
  NOR2_X1 U16902 ( .A1(net749636), .A2(net765546), .ZN(net714842) );
  AND2_X1 U16903 ( .A1(net715146), .A2(net713607), .ZN(net758037) );
  NOR2_X1 U16904 ( .A1(net715146), .A2(net713607), .ZN(net714602) );
  NAND2_X1 U16905 ( .A1(net714008), .A2(net741987), .ZN(net713467) );
  NOR2_X1 U16906 ( .A1(net725077), .A2(net745681), .ZN(net745679) );
  INV_X1 U16907 ( .A(net725077), .ZN(net749442) );
  NAND2_X1 U16908 ( .A1(net714002), .A2(net714007), .ZN(net731199) );
  NAND3_X1 U16909 ( .A1(net717591), .A2(net742326), .A3(net730300), .ZN(
        net738443) );
  NAND3_X1 U16910 ( .A1(net714612), .A2(net767213), .A3(net714611), .ZN(
        net726959) );
  OAI21_X1 U16911 ( .B1(net714611), .B2(net750290), .A(net767213), .ZN(
        net728159) );
  NAND2_X1 U16912 ( .A1(net750290), .A2(net767213), .ZN(net726961) );
  CLKBUF_X1 U16913 ( .A(net718140), .Z(net786867) );
  AND2_X2 U16914 ( .A1(net749307), .A2(net718140), .ZN(net742326) );
  INV_X1 U16915 ( .A(net714119), .ZN(net714122) );
  AND2_X1 U16916 ( .A1(net714845), .A2(net714119), .ZN(net749307) );
  INV_X1 U16917 ( .A(net714842), .ZN(net746753) );
  INV_X1 U16918 ( .A(net717967), .ZN(net716249) );
  AOI21_X1 U16919 ( .B1(n6461), .B2(net712797), .A(net712810), .ZN(n22866) );
  NAND2_X1 U16920 ( .A1(net712795), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [20]), .ZN(net712797) );
  NOR3_X1 U16921 ( .A1(net749439), .A2(n6461), .A3(net780298), .ZN(net712810)
         );
  CLKBUF_X3 U16922 ( .A(net717950), .Z(net716341) );
  XNOR2_X1 U16923 ( .A(net745672), .B(net745684), .ZN(net749239) );
  NOR2_X1 U16924 ( .A1(net741456), .A2(net366451), .ZN(net712459) );
  AOI21_X1 U16925 ( .B1(net712855), .B2(net732762), .A(net732750), .ZN(
        net713973) );
  AOI22_X1 U16926 ( .A1(net713873), .A2(net767211), .B1(net713979), .B2(
        net713874), .ZN(net713974) );
  NAND2_X1 U16927 ( .A1(net713978), .A2(net713779), .ZN(net713975) );
  NAND2_X1 U16928 ( .A1(net713869), .A2(net713785), .ZN(net713976) );
  NOR2_X1 U16929 ( .A1(n6461), .A2(net749434), .ZN(net780360) );
  OAI21_X1 U16930 ( .B1(net712795), .B2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [20]), .A(net712797), .ZN(net712794) );
  OAI21_X1 U16931 ( .B1(net712810), .B2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [22]), .A(net712812), .ZN(net712809) );
  OR2_X1 U16932 ( .A1(net713909), .A2(net734493), .ZN(net780215) );
  NAND2_X1 U16933 ( .A1(net741999), .A2(n22685), .ZN(n23193) );
  INV_X1 U16934 ( .A(net787514), .ZN(net787526) );
  INV_X1 U16935 ( .A(net787514), .ZN(net787528) );
  NOR2_X1 U16936 ( .A1(net712812), .A2(n6462), .ZN(n26570) );
  AND2_X1 U16937 ( .A1(net741999), .A2(s_IFID_IR[23]), .ZN(n22867) );
  BUF_X2 U16938 ( .A(net713853), .Z(net718405) );
  OR2_X1 U16939 ( .A1(net716341), .A2(n23467), .ZN(n26712) );
  AND3_X2 U16940 ( .A1(n23763), .A2(n24138), .A3(n23764), .ZN(n23949) );
  OAI21_X1 U16941 ( .B1(n26129), .B2(n26128), .A(n26127), .ZN(n22868) );
  INV_X1 U16942 ( .A(net713564), .ZN(net786856) );
  INV_X1 U16943 ( .A(net713564), .ZN(net713868) );
  BUF_X2 U16944 ( .A(net713868), .Z(net755699) );
  CLKBUF_X1 U16945 ( .A(n24136), .Z(n22869) );
  MUX2_X1 U16946 ( .A(\core_inst/EXMEM_NPC/DFF_13/N3 ), .B(n26077), .S(
        net716237), .Z(n26042) );
  BUF_X1 U16947 ( .A(n25766), .Z(n22870) );
  NAND2_X1 U16948 ( .A1(n24320), .A2(n25319), .ZN(n25416) );
  BUF_X1 U16949 ( .A(n24360), .Z(n23993) );
  CLKBUF_X3 U16950 ( .A(net717844), .Z(net742092) );
  BUF_X2 U16951 ( .A(net717844), .Z(net742339) );
  INV_X1 U16952 ( .A(net718340), .ZN(net786841) );
  BUF_X1 U16953 ( .A(net749922), .Z(net786837) );
  NOR2_X1 U16954 ( .A1(n23604), .A2(n24192), .ZN(n22871) );
  OR2_X1 U16955 ( .A1(net89524), .A2(net715769), .ZN(n22872) );
  OR2_X1 U16956 ( .A1(n22872), .A2(net742011), .ZN(n23941) );
  CLKBUF_X2 U16957 ( .A(net718372), .Z(net749387) );
  OAI222_X4 U16958 ( .A1(n26031), .A2(n25909), .B1(net762754), .B2(n24577), 
        .C1(net717055), .C2(net713701), .ZN(n25912) );
  INV_X1 U16959 ( .A(net762579), .ZN(net718133) );
  INV_X1 U16960 ( .A(net714631), .ZN(net786824) );
  NOR2_X1 U16961 ( .A1(n23006), .A2(n23007), .ZN(n22873) );
  AND3_X1 U16962 ( .A1(n22835), .A2(net749338), .A3(net749905), .ZN(net749428)
         );
  OR2_X1 U16963 ( .A1(net716341), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_g[2] ), .ZN(n26719) );
  INV_X1 U16964 ( .A(net714248), .ZN(net765428) );
  OAI21_X1 U16965 ( .B1(n24525), .B2(net714689), .A(n23642), .ZN(n25791) );
  INV_X1 U16966 ( .A(net796014), .ZN(net765429) );
  OAI222_X1 U16967 ( .A1(net755631), .A2(net713683), .B1(n24572), .B2(n24548), 
        .C1(net713707), .C2(net714689), .ZN(n23540) );
  NOR2_X1 U16968 ( .A1(net796014), .A2(net742243), .ZN(n22975) );
  NAND2_X1 U16969 ( .A1(net749886), .A2(n24341), .ZN(net715014) );
  NAND2_X1 U16970 ( .A1(net749886), .A2(net713614), .ZN(n25884) );
  CLKBUF_X1 U16971 ( .A(net715014), .Z(net749839) );
  NAND3_X1 U16972 ( .A1(n26043), .A2(net714275), .A3(n22875), .ZN(n23707) );
  NAND2_X1 U16973 ( .A1(n26148), .A2(net750019), .ZN(n22875) );
  NAND4_X1 U16974 ( .A1(n22875), .A2(n26044), .A3(n26045), .A4(n26043), .ZN(
        n22880) );
  NAND2_X1 U16975 ( .A1(n22879), .A2(net715555), .ZN(n22876) );
  OAI22_X1 U16976 ( .A1(net767209), .A2(n22876), .B1(n22881), .B2(net714267), 
        .ZN(n22878) );
  OAI222_X1 U16977 ( .A1(n26174), .A2(net767209), .B1(n26055), .B2(net748269), 
        .C1(n22876), .C2(net767210), .ZN(n25869) );
  NAND2_X1 U16978 ( .A1(n22876), .A2(net713733), .ZN(n26178) );
  OAI222_X1 U16979 ( .A1(n26173), .A2(net767209), .B1(net713154), .B2(n25796), 
        .C1(net714267), .C2(n22876), .ZN(n25805) );
  AND2_X2 U16980 ( .A1(n24331), .A2(n25371), .ZN(n22877) );
  AOI22_X1 U16981 ( .A1(n25797), .A2(net713775), .B1(n22877), .B2(net714275), 
        .ZN(n25803) );
  NAND2_X1 U16982 ( .A1(n22877), .A2(net767208), .ZN(n24398) );
  NAND2_X1 U16983 ( .A1(n22877), .A2(net714306), .ZN(n22899) );
  NOR2_X1 U16984 ( .A1(n22878), .A2(n25765), .ZN(n22932) );
  BUF_X1 U16985 ( .A(n22878), .Z(n23026) );
  CLKBUF_X1 U16986 ( .A(net731393), .Z(net734607) );
  INV_X1 U16987 ( .A(net795993), .ZN(net716369) );
  INV_X1 U16988 ( .A(net742612), .ZN(net716367) );
  NOR2_X1 U16989 ( .A1(net765428), .A2(net750255), .ZN(net742247) );
  AOI22_X1 U16990 ( .A1(n22880), .A2(net749534), .B1(net749500), .B2(n24539), 
        .ZN(n22879) );
  AND2_X1 U16991 ( .A1(n25774), .A2(n25761), .ZN(n22882) );
  NAND3_X1 U16992 ( .A1(n24259), .A2(n25762), .A3(n22882), .ZN(n22881) );
  OAI22_X1 U16993 ( .A1(net750203), .A2(n24279), .B1(n25600), .B2(net713564), 
        .ZN(net786066) );
  OR2_X1 U16994 ( .A1(net713990), .A2(n24547), .ZN(n22883) );
  AND2_X1 U16995 ( .A1(n22883), .A2(n25774), .ZN(n25371) );
  CLKBUF_X1 U16996 ( .A(n25447), .Z(n22901) );
  MUX2_X1 U16997 ( .A(net713892), .B(n26136), .S(n24318), .Z(n22892) );
  OAI22_X1 U16998 ( .A1(net748269), .A2(net750287), .B1(net762754), .B2(
        net750274), .ZN(n22887) );
  OAI222_X1 U16999 ( .A1(net728314), .A2(net762661), .B1(net717055), .B2(
        n24358), .C1(net717074), .C2(net742483), .ZN(n22886) );
  INV_X1 U17000 ( .A(n26037), .ZN(n22896) );
  INV_X1 U17001 ( .A(n26036), .ZN(n22895) );
  NAND2_X1 U17002 ( .A1(n22901), .A2(n24308), .ZN(n22897) );
  NOR2_X1 U17003 ( .A1(n26038), .A2(n22892), .ZN(n22891) );
  MUX2_X1 U17004 ( .A(net713728), .B(net717087), .S(n24318), .Z(n22890) );
  OAI21_X1 U17005 ( .B1(n22886), .B2(n22887), .A(net713775), .ZN(n22885) );
  OAI211_X1 U17006 ( .C1(n24332), .C2(n22895), .A(n24308), .B(n22896), .ZN(
        n22894) );
  NAND3_X1 U17007 ( .A1(n22897), .A2(n26037), .A3(n26036), .ZN(n22893) );
  NAND2_X1 U17008 ( .A1(n24545), .A2(net749710), .ZN(n22900) );
  MUX2_X1 U17009 ( .A(n22890), .B(n22891), .S(net780543), .Z(n22888) );
  NAND2_X1 U17010 ( .A1(n26039), .A2(net714275), .ZN(n22889) );
  OAI21_X1 U17011 ( .B1(n26040), .B2(net714267), .A(n22885), .ZN(n22884) );
  AND3_X1 U17012 ( .A1(n22893), .A2(net717091), .A3(n22894), .ZN(n22898) );
  AND4_X1 U17013 ( .A1(n22899), .A2(n22889), .A3(n22888), .A4(n22900), .ZN(
        net749219) );
  NOR2_X1 U17014 ( .A1(n22898), .A2(n22884), .ZN(net717684) );
  INV_X1 U17015 ( .A(n25600), .ZN(n22905) );
  NAND2_X1 U17016 ( .A1(n22905), .A2(n22980), .ZN(n22904) );
  NOR2_X1 U17017 ( .A1(n25789), .A2(n24274), .ZN(n22902) );
  AOI211_X1 U17018 ( .C1(net767206), .C2(net717463), .A(n22902), .B(n22903), 
        .ZN(n25784) );
  NAND2_X1 U17019 ( .A1(n22904), .A2(n25884), .ZN(n22903) );
  NAND3_X1 U17020 ( .A1(n26158), .A2(n26156), .A3(n26155), .ZN(n22908) );
  NAND3_X1 U17021 ( .A1(n26154), .A2(net767211), .A3(n26157), .ZN(n22907) );
  NAND2_X1 U17022 ( .A1(n25784), .A2(n25783), .ZN(n22906) );
  OAI22_X1 U17023 ( .A1(n22906), .A2(net713897), .B1(n22907), .B2(n22908), 
        .ZN(n26409) );
  INV_X1 U17024 ( .A(n26566), .ZN(n22924) );
  NAND3_X1 U17025 ( .A1(n25366), .A2(n26566), .A3(net713751), .ZN(n22925) );
  INV_X1 U17026 ( .A(n25875), .ZN(n22920) );
  BUF_X1 U17027 ( .A(n25405), .Z(n22935) );
  NOR3_X1 U17028 ( .A1(n25875), .A2(net749289), .A3(n23023), .ZN(n22923) );
  NOR3_X1 U17029 ( .A1(n22924), .A2(net713863), .A3(n26565), .ZN(n22922) );
  OAI21_X1 U17030 ( .B1(n26560), .B2(n25875), .A(n22925), .ZN(n22921) );
  NOR2_X1 U17031 ( .A1(n26563), .A2(net713863), .ZN(n22926) );
  AOI21_X1 U17032 ( .B1(net713951), .B2(net713949), .A(n26409), .ZN(n22931) );
  NOR2_X1 U17033 ( .A1(n24234), .A2(n24399), .ZN(n22933) );
  NAND2_X1 U17034 ( .A1(n22935), .A2(n22920), .ZN(n22919) );
  NOR3_X1 U17035 ( .A1(n22921), .A2(n22922), .A3(n22923), .ZN(n22918) );
  AND4_X1 U17036 ( .A1(n22926), .A2(net749289), .A3(n26566), .A4(net714934), 
        .ZN(n22934) );
  OAI211_X1 U17037 ( .C1(n25769), .C2(n25768), .A(n22932), .B(n25767), .ZN(
        n13082) );
  NAND3_X1 U17038 ( .A1(n22931), .A2(n26406), .A3(n26407), .ZN(n22930) );
  NAND3_X1 U17039 ( .A1(n24397), .A2(n24398), .A3(n22933), .ZN(n22911) );
  NOR2_X1 U17040 ( .A1(n25933), .A2(n25338), .ZN(n22912) );
  NOR2_X1 U17041 ( .A1(n25415), .A2(n26533), .ZN(n22914) );
  NAND3_X1 U17042 ( .A1(net713448), .A2(net717091), .A3(net714105), .ZN(n22913) );
  OAI211_X1 U17043 ( .C1(net717091), .C2(n26567), .A(n22918), .B(n22919), .ZN(
        n22917) );
  NOR3_X1 U17044 ( .A1(n23397), .A2(n23023), .A3(n25875), .ZN(n22916) );
  AND2_X1 U17045 ( .A1(n25502), .A2(n22934), .ZN(n22915) );
  AOI21_X1 U17046 ( .B1(n24382), .B2(net717091), .A(n24383), .ZN(n22909) );
  AOI21_X1 U17047 ( .B1(n24235), .B2(net717091), .A(n24236), .ZN(n22910) );
  NAND3_X1 U17048 ( .A1(net728481), .A2(net714335), .A3(net717091), .ZN(n22927) );
  NOR2_X1 U17049 ( .A1(n13082), .A2(n26607), .ZN(n22929) );
  NOR3_X1 U17050 ( .A1(n25512), .A2(n22911), .A3(n22930), .ZN(n22928) );
  OR2_X1 U17051 ( .A1(n26529), .A2(n25383), .ZN(net740704) );
  OAI211_X1 U17052 ( .C1(net712494), .C2(net713154), .A(net712493), .B(n22912), 
        .ZN(net714732) );
  NAND3_X1 U17053 ( .A1(n22913), .A2(n26580), .A3(n22914), .ZN(net714622) );
  NOR3_X1 U17054 ( .A1(n22915), .A2(n22916), .A3(n22917), .ZN(net714911) );
  NAND4_X1 U17055 ( .A1(n26724), .A2(n22927), .A3(n22910), .A4(n22909), .ZN(
        net714910) );
  NAND4_X1 U17056 ( .A1(n22928), .A2(n22929), .A3(n26726), .A4(n26606), .ZN(
        net714909) );
  NOR3_X1 U17057 ( .A1(net712838), .A2(n6402), .A3(net780340), .ZN(net712886)
         );
  NOR2_X2 U17058 ( .A1(n26576), .A2(n6460), .ZN(n26575) );
  AND2_X2 U17059 ( .A1(net780532), .A2(net755005), .ZN(n22936) );
  AND2_X2 U17060 ( .A1(net780532), .A2(net755005), .ZN(n24260) );
  INV_X1 U17061 ( .A(n26707), .ZN(n22938) );
  NOR2_X1 U17062 ( .A1(net796143), .A2(n22674), .ZN(
        \core_inst/EXMEM_RF_ADDR_DEST/DFF_0/N3 ) );
  AND2_X1 U17063 ( .A1(net742649), .A2(n25588), .ZN(n22939) );
  NOR2_X1 U17064 ( .A1(net796143), .A2(n23297), .ZN(n23984) );
  AND2_X1 U17065 ( .A1(net716255), .A2(n18059), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_1/N3 ) );
  AND2_X1 U17066 ( .A1(net716267), .A2(n22942), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_5/N3 ) );
  AND2_X1 U17067 ( .A1(net741999), .A2(n22944), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_15/N3 ) );
  AND2_X1 U17068 ( .A1(net716259), .A2(s_IFID_IR[20]), .ZN(n22945) );
  INV_X1 U17069 ( .A(net716265), .ZN(net785270) );
  BUF_X1 U17070 ( .A(n26561), .Z(n23023) );
  INV_X1 U17071 ( .A(net716341), .ZN(net742648) );
  INV_X1 U17072 ( .A(net716341), .ZN(net716267) );
  INV_X1 U17073 ( .A(net716337), .ZN(net716253) );
  MUX2_X1 U17074 ( .A(n790), .B(n26101), .S(net787528), .Z(net713777) );
  AND2_X1 U17075 ( .A1(net716253), .A2(n22946), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_13/N3 ) );
  AND2_X1 U17076 ( .A1(net716247), .A2(n23938), .ZN(n22947) );
  INV_X1 U17077 ( .A(net742576), .ZN(net785239) );
  BUF_X1 U17078 ( .A(n25402), .Z(n22948) );
  NAND2_X1 U17079 ( .A1(n23011), .A2(net740674), .ZN(n22949) );
  BUF_X2 U17080 ( .A(net713853), .Z(net785220) );
  BUF_X2 U17081 ( .A(net713853), .Z(net785219) );
  NAND2_X1 U17082 ( .A1(n23934), .A2(net715700), .ZN(net742257) );
  INV_X1 U17083 ( .A(net742257), .ZN(net715592) );
  INV_X1 U17084 ( .A(net796159), .ZN(net714943) );
  BUF_X1 U17085 ( .A(net796159), .Z(net742017) );
  INV_X1 U17086 ( .A(net796159), .ZN(net749495) );
  INV_X1 U17087 ( .A(net713844), .ZN(net780582) );
  CLKBUF_X1 U17088 ( .A(net713844), .Z(net780566) );
  AND2_X1 U17089 ( .A1(net713844), .A2(n17667), .ZN(n23449) );
  INV_X1 U17090 ( .A(net713844), .ZN(net765629) );
  INV_X1 U17091 ( .A(net713844), .ZN(net715058) );
  NAND2_X1 U17092 ( .A1(net713844), .A2(n25334), .ZN(n25754) );
  INV_X1 U17093 ( .A(net713844), .ZN(net749926) );
  INV_X1 U17094 ( .A(net713844), .ZN(net717615) );
  CLKBUF_X1 U17095 ( .A(net713844), .Z(net742331) );
  CLKBUF_X1 U17096 ( .A(net713844), .Z(net749806) );
  INV_X1 U17097 ( .A(net713844), .ZN(net742037) );
  CLKBUF_X1 U17098 ( .A(net741980), .Z(net780522) );
  NOR2_X1 U17099 ( .A1(net741980), .A2(n25384), .ZN(n25585) );
  OR2_X2 U17100 ( .A1(net717845), .A2(net732423), .ZN(net717543) );
  CLKBUF_X1 U17101 ( .A(net732423), .Z(net717570) );
  INV_X1 U17102 ( .A(net749316), .ZN(net717844) );
  INV_X1 U17103 ( .A(net749316), .ZN(net717845) );
  XNOR2_X1 U17104 ( .A(net749316), .B(net716215), .ZN(n25793) );
  AND2_X2 U17105 ( .A1(net717844), .A2(net755214), .ZN(n22950) );
  AND2_X1 U17106 ( .A1(net717844), .A2(net755214), .ZN(n25420) );
  NAND3_X1 U17107 ( .A1(net717844), .A2(n25577), .A3(n24567), .ZN(n25389) );
  NOR2_X1 U17108 ( .A1(net717844), .A2(n24567), .ZN(n26022) );
  BUF_X1 U17109 ( .A(net714248), .Z(net750057) );
  INV_X1 U17110 ( .A(net714248), .ZN(net749273) );
  INV_X1 U17111 ( .A(net714248), .ZN(net714689) );
  NOR2_X1 U17112 ( .A1(net765428), .A2(n26193), .ZN(n23323) );
  NAND3_X1 U17113 ( .A1(n22950), .A2(net715313), .A3(n24566), .ZN(net713853)
         );
  AOI22_X1 U17114 ( .A1(n23346), .A2(n22950), .B1(net750025), .B2(net718391), 
        .ZN(n25775) );
  AOI22_X1 U17115 ( .A1(n23360), .A2(n22950), .B1(net750158), .B2(n24345), 
        .ZN(n25771) );
  AOI22_X1 U17116 ( .A1(net749525), .A2(n22950), .B1(net749306), .B2(net750057), .ZN(n23460) );
  AOI211_X1 U17117 ( .C1(n22950), .C2(net755238), .A(net750255), .B(net713882), 
        .ZN(n25432) );
  AOI22_X1 U17118 ( .A1(net742506), .A2(n22950), .B1(net750238), .B2(net750057), .ZN(n25899) );
  NAND2_X1 U17119 ( .A1(n22950), .A2(net755241), .ZN(n25426) );
  OAI222_X1 U17120 ( .A1(n25578), .A2(net718405), .B1(net713907), .B2(
        net713868), .C1(net750278), .C2(net742259), .ZN(net714389) );
  OAI22_X1 U17121 ( .A1(net713907), .A2(n24358), .B1(net718405), .B2(net742271), .ZN(n23000) );
  OAI222_X1 U17122 ( .A1(net713907), .A2(net742087), .B1(net785220), .B2(
        net786856), .C1(n24303), .C2(net731327), .ZN(net714431) );
  OAI222_X1 U17123 ( .A1(n25578), .A2(net713907), .B1(net785219), .B2(
        net713905), .C1(net717055), .C2(net749454), .ZN(n25930) );
  INV_X1 U17124 ( .A(net785219), .ZN(net713748) );
  OAI222_X1 U17125 ( .A1(net718405), .A2(n24269), .B1(n24310), .B2(net749823), 
        .C1(net713907), .C2(net742483), .ZN(n25880) );
  OAI22_X1 U17126 ( .A1(n24303), .A2(net742271), .B1(net718405), .B2(net748269), .ZN(n24394) );
  NOR2_X1 U17127 ( .A1(net785220), .A2(net742087), .ZN(n24409) );
  OAI222_X1 U17128 ( .A1(net762754), .A2(net713701), .B1(n26031), .B2(n24539), 
        .C1(net785219), .C2(net742483), .ZN(n26032) );
  AND3_X1 U17129 ( .A1(n24560), .A2(n24310), .A3(net718405), .ZN(net712469) );
  OAI22_X1 U17130 ( .A1(net713907), .A2(net755238), .B1(net785220), .B2(
        net749823), .ZN(n25913) );
  NAND4_X1 U17131 ( .A1(net713907), .A2(n24270), .A3(net755683), .A4(net785219), .ZN(n26008) );
  OAI22_X1 U17132 ( .A1(net785220), .A2(net742259), .B1(n26031), .B2(n24341), 
        .ZN(n25948) );
  OAI211_X1 U17133 ( .C1(net780556), .C2(n24274), .A(n22954), .B(n22955), .ZN(
        n22951) );
  NOR2_X1 U17134 ( .A1(n22952), .A2(n22951), .ZN(n24331) );
  NAND2_X1 U17135 ( .A1(net750024), .A2(n25586), .ZN(n22953) );
  OAI21_X1 U17136 ( .B1(net749685), .B2(n25789), .A(n22953), .ZN(n22952) );
  AOI21_X1 U17137 ( .B1(n24272), .B2(net717875), .A(net784601), .ZN(n22954) );
  NAND2_X1 U17138 ( .A1(n24401), .A2(n24341), .ZN(n22955) );
  MUX2_X1 U17139 ( .A(net713728), .B(net713770), .S(n26199), .Z(n22958) );
  MUX2_X1 U17140 ( .A(net713726), .B(n25662), .S(n26199), .Z(n22957) );
  NAND2_X1 U17141 ( .A1(n26023), .A2(net742339), .ZN(n22964) );
  NOR2_X1 U17142 ( .A1(n25443), .A2(net748274), .ZN(n22962) );
  INV_X1 U17143 ( .A(n25663), .ZN(n22961) );
  MUX2_X1 U17144 ( .A(n22957), .B(n22958), .S(net750019), .Z(n22956) );
  NAND4_X1 U17145 ( .A1(n22964), .A2(n25451), .A3(net767211), .A4(n24536), 
        .ZN(n22963) );
  AOI21_X1 U17146 ( .B1(n24550), .B2(net749685), .A(n22962), .ZN(n22960) );
  AOI22_X1 U17147 ( .A1(n25402), .A2(net714394), .B1(n22961), .B2(n24525), 
        .ZN(n22959) );
  NOR2_X1 U17148 ( .A1(net714382), .A2(n24030), .ZN(net714380) );
  NAND2_X1 U17149 ( .A1(n22963), .A2(n22956), .ZN(net714379) );
  OAI222_X1 U17150 ( .A1(net717056), .A2(net718391), .B1(net748275), .B2(
        net750019), .C1(net717059), .C2(net718380), .ZN(net714388) );
  OAI222_X1 U17151 ( .A1(n24291), .A2(net713773), .B1(net717053), .B2(
        net742508), .C1(net713851), .C2(net713905), .ZN(net714387) );
  NAND2_X1 U17152 ( .A1(n22960), .A2(n22959), .ZN(net714386) );
  NOR2_X2 U17153 ( .A1(n25411), .A2(n22965), .ZN(n25923) );
  NOR2_X2 U17154 ( .A1(n26063), .A2(net784220), .ZN(n22965) );
  INV_X2 U17155 ( .A(net734022), .ZN(net784220) );
  NOR2_X1 U17156 ( .A1(net715365), .A2(n24267), .ZN(n22966) );
  NOR2_X1 U17157 ( .A1(n22966), .A2(n23029), .ZN(n23019) );
  NOR2_X1 U17158 ( .A1(n22966), .A2(n26062), .ZN(n23732) );
  NAND2_X1 U17159 ( .A1(n22975), .A2(n24577), .ZN(net715021) );
  NAND3_X1 U17160 ( .A1(net715019), .A2(net715020), .A3(net715021), .ZN(n24246) );
  NAND4_X1 U17161 ( .A1(net731685), .A2(net715018), .A3(net715019), .A4(
        net715020), .ZN(n23766) );
  INV_X1 U17162 ( .A(net716339), .ZN(net716265) );
  OR2_X1 U17163 ( .A1(net796200), .A2(n24527), .ZN(n26720) );
  OR3_X1 U17164 ( .A1(net765730), .A2(n25622), .A3(net716339), .ZN(n24427) );
  INV_X1 U17165 ( .A(net716339), .ZN(net765341) );
  INV_X1 U17166 ( .A(net716339), .ZN(net716247) );
  INV_X1 U17167 ( .A(net716339), .ZN(net716257) );
  INV_X1 U17168 ( .A(net765340), .ZN(n15091) );
  BUF_X1 U17169 ( .A(n15091), .Z(net742612) );
  INV_X1 U17170 ( .A(net795993), .ZN(net716377) );
  NAND2_X1 U17171 ( .A1(net716385), .A2(s_IFID_IR[17]), .ZN(n26569) );
  AND2_X1 U17172 ( .A1(net742576), .A2(n17722), .ZN(
        \core_inst/IDEX_NPC/DFF_27/N3 ) );
  NOR2_X1 U17173 ( .A1(net716367), .A2(n24334), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_4/N3 ) );
  NOR2_X1 U17174 ( .A1(net796137), .A2(n5595), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_24/N3 ) );
  NOR2_X1 U17175 ( .A1(net716333), .A2(n5618), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_7/N3 ) );
  INV_X1 U17176 ( .A(net717952), .ZN(net742084) );
  OAI211_X1 U17177 ( .C1(n25747), .C2(n24316), .A(n24135), .B(
        \cu_inst/FW_UNIT/ITD_EXMEM/N14 ), .ZN(net715799) );
  XNOR2_X1 U17178 ( .A(n1668), .B(n1641), .ZN(n22971) );
  XNOR2_X1 U17179 ( .A(net718087), .B(n5181), .ZN(n22970) );
  XOR2_X1 U17180 ( .A(net742084), .B(n5607), .Z(n22972) );
  XOR2_X1 U17181 ( .A(net717830), .B(\core_inst/MEMWB_IR/DFF_15/N3 ), .Z(
        n22973) );
  XNOR2_X1 U17182 ( .A(net718083), .B(n1637), .ZN(n22974) );
  NAND2_X1 U17183 ( .A1(n22970), .A2(n22971), .ZN(n22969) );
  NAND3_X1 U17184 ( .A1(n22974), .A2(n22973), .A3(n22972), .ZN(n22968) );
  INV_X1 U17185 ( .A(net715692), .ZN(net715721) );
  NOR2_X1 U17186 ( .A1(n22968), .A2(n22969), .ZN(n22967) );
  NAND3_X1 U17187 ( .A1(n22967), .A2(n25750), .A3(net715721), .ZN(n23947) );
  OR2_X1 U17188 ( .A1(net717543), .A2(net749698), .ZN(n24267) );
  INV_X1 U17189 ( .A(net715284), .ZN(net715365) );
  NAND2_X1 U17190 ( .A1(n22979), .A2(n25940), .ZN(n22976) );
  NOR2_X1 U17191 ( .A1(n22976), .A2(net718103), .ZN(net714706) );
  AND2_X1 U17192 ( .A1(n22979), .A2(n25940), .ZN(n23888) );
  OAI22_X1 U17193 ( .A1(net715420), .A2(n4401), .B1(n1710), .B2(net718154), 
        .ZN(n22978) );
  OAI22_X1 U17194 ( .A1(n23266), .A2(net715421), .B1(net717719), .B2(n4400), 
        .ZN(n22977) );
  NOR2_X1 U17195 ( .A1(n22977), .A2(n22978), .ZN(net714077) );
  MUX2_X2 U17196 ( .A(n1064), .B(net714077), .S(net787526), .Z(n26149) );
  NAND2_X1 U17197 ( .A1(n25840), .A2(n24555), .ZN(n24288) );
  NAND2_X1 U17198 ( .A1(n24288), .A2(n25936), .ZN(n22979) );
  XOR2_X1 U17199 ( .A(n24302), .B(n22980), .Z(net783467) );
  NOR2_X1 U17200 ( .A1(n23920), .A2(net714287), .ZN(n22981) );
  AOI21_X1 U17201 ( .B1(n22981), .B2(net783470), .A(n22982), .ZN(net783466) );
  INV_X1 U17202 ( .A(n22844), .ZN(net783470) );
  OAI21_X1 U17203 ( .B1(n23920), .B2(net741987), .A(n24361), .ZN(n22982) );
  NAND2_X1 U17204 ( .A1(n24298), .A2(net749375), .ZN(n25766) );
  NOR2_X1 U17205 ( .A1(n25766), .A2(net749698), .ZN(n25779) );
  NAND3_X1 U17206 ( .A1(n25779), .A2(net718367), .A3(net717511), .ZN(net713866) );
  XNOR2_X1 U17207 ( .A(net786821), .B(net713711), .ZN(n23832) );
  INV_X1 U17208 ( .A(net717967), .ZN(net742368) );
  NAND2_X1 U17209 ( .A1(net716249), .A2(s_IFID_IR[18]), .ZN(n23953) );
  NAND3_X1 U17210 ( .A1(net716249), .A2(net717049), .A3(n26603), .ZN(n25537)
         );
  AND2_X1 U17211 ( .A1(net716259), .A2(n17940), .ZN(
        \core_inst/IDEX_NPC/DFF_6/N3 ) );
  AND2_X1 U17212 ( .A1(net785255), .A2(n17785), .ZN(
        \core_inst/IDEX_NPC/DFF_18/N3 ) );
  OAI21_X1 U17213 ( .B1(n26740), .B2(net760161), .A(n26582), .ZN(
        \core_inst/IF_stage/PROGRAM_COUNTER/DFF_0/N3 ) );
  AND2_X1 U17214 ( .A1(net741999), .A2(n25446), .ZN(n23992) );
  AND2_X1 U17215 ( .A1(net742649), .A2(n26257), .ZN(n23991) );
  NOR2_X2 U17216 ( .A1(n25872), .A2(net786856), .ZN(n26129) );
  OAI21_X1 U17217 ( .B1(n26129), .B2(n26128), .A(n26127), .ZN(n24096) );
  OAI21_X1 U17218 ( .B1(n25366), .B2(n26130), .A(n24096), .ZN(n24309) );
  NAND2_X1 U17219 ( .A1(n24309), .A2(net718400), .ZN(net731060) );
  NAND3_X1 U17220 ( .A1(net782764), .A2(n22984), .A3(n22983), .ZN(n25988) );
  NAND2_X1 U17221 ( .A1(net713614), .A2(n24190), .ZN(n22984) );
  AOI22_X1 U17222 ( .A1(net714251), .A2(net742242), .B1(n24577), .B2(n22673), 
        .ZN(n22983) );
  MUX2_X1 U17223 ( .A(n25988), .B(n25920), .S(net750176), .Z(net713894) );
  NAND2_X1 U17224 ( .A1(net714657), .A2(net714309), .ZN(n25414) );
  OAI22_X1 U17225 ( .A1(net717059), .A2(net718391), .B1(net718406), .B2(
        net748274), .ZN(n22987) );
  INV_X1 U17226 ( .A(net717053), .ZN(net727843) );
  NOR2_X1 U17227 ( .A1(net717056), .A2(net731327), .ZN(n22991) );
  OAI22_X1 U17228 ( .A1(n24338), .A2(net742506), .B1(net755241), .B2(n25663), 
        .ZN(n22990) );
  NAND2_X1 U17229 ( .A1(n24203), .A2(net734022), .ZN(n22986) );
  INV_X1 U17230 ( .A(n22987), .ZN(n22985) );
  NAND2_X1 U17231 ( .A1(net727843), .A2(net714494), .ZN(n22989) );
  NOR2_X1 U17232 ( .A1(n22990), .A2(n22991), .ZN(n22988) );
  INV_X1 U17233 ( .A(net713874), .ZN(net727832) );
  OAI211_X1 U17234 ( .C1(n24310), .C2(net755699), .A(n22985), .B(n22986), .ZN(
        net727834) );
  OAI211_X1 U17235 ( .C1(n25599), .C2(net767206), .A(n22988), .B(n22989), .ZN(
        net727833) );
  NOR2_X1 U17236 ( .A1(n26135), .A2(net727832), .ZN(net727831) );
  OAI22_X1 U17237 ( .A1(net713882), .A2(n25448), .B1(net749454), .B2(net713767), .ZN(net727830) );
  OAI22_X1 U17238 ( .A1(n24303), .A2(n24269), .B1(n24560), .B2(net767207), 
        .ZN(n23005) );
  NAND2_X1 U17239 ( .A1(net712466), .A2(net780543), .ZN(n23004) );
  INV_X1 U17240 ( .A(n23005), .ZN(n23003) );
  INV_X1 U17241 ( .A(n25969), .ZN(n22996) );
  NAND3_X1 U17242 ( .A1(n25414), .A2(net767203), .A3(n25968), .ZN(n22995) );
  OAI22_X1 U17243 ( .A1(net762754), .A2(net717875), .B1(net713701), .B2(n26031), .ZN(n22999) );
  OAI22_X1 U17244 ( .A1(net749387), .A2(net717074), .B1(n24357), .B2(net749525), .ZN(n22998) );
  OAI22_X1 U17245 ( .A1(net749822), .A2(net717055), .B1(n24270), .B2(net748269), .ZN(n22997) );
  NAND3_X1 U17246 ( .A1(n25414), .A2(n23003), .A3(n23004), .ZN(n23001) );
  NAND2_X1 U17247 ( .A1(n25968), .A2(n25969), .ZN(n23002) );
  NOR3_X1 U17248 ( .A1(n22995), .A2(n22996), .A3(n25970), .ZN(n22994) );
  NOR4_X1 U17249 ( .A1(n22997), .A2(n22998), .A3(n22999), .A4(n23000), .ZN(
        n22993) );
  NOR3_X1 U17250 ( .A1(n25970), .A2(n23002), .A3(n23001), .ZN(n22992) );
  AOI21_X1 U17251 ( .B1(n22992), .B2(n22993), .A(n22994), .ZN(n25415) );
  NAND3_X1 U17252 ( .A1(net796122), .A2(net366126), .A3(net749369), .ZN(n23008) );
  OR2_X1 U17253 ( .A1(net749951), .A2(net715460), .ZN(n23010) );
  NAND3_X1 U17254 ( .A1(net717876), .A2(net749664), .A3(n14764), .ZN(n23009)
         );
  OAI21_X1 U17255 ( .B1(n23010), .B2(n1690), .A(n23008), .ZN(n23007) );
  OAI21_X1 U17256 ( .B1(net717718), .B2(n4418), .A(n23009), .ZN(n23006) );
  NOR2_X1 U17257 ( .A1(n23006), .A2(n23007), .ZN(n26099) );
  NAND2_X1 U17258 ( .A1(n26099), .A2(net787512), .ZN(n23011) );
  NAND2_X1 U17259 ( .A1(n23011), .A2(net740674), .ZN(n26185) );
  NAND2_X1 U17260 ( .A1(net750228), .A2(n24206), .ZN(n23012) );
  NAND2_X1 U17261 ( .A1(n22949), .A2(net750255), .ZN(n23014) );
  NAND3_X1 U17262 ( .A1(n24341), .A2(n24566), .A3(net717570), .ZN(n23013) );
  NAND4_X1 U17263 ( .A1(n24558), .A2(n23013), .A3(n23014), .A4(n23012), .ZN(
        n25920) );
  NAND2_X1 U17264 ( .A1(n25920), .A2(net742092), .ZN(n26026) );
  NAND2_X1 U17265 ( .A1(net749317), .A2(net713701), .ZN(net781609) );
  AND2_X1 U17266 ( .A1(n26024), .A2(n26027), .ZN(n23015) );
  NAND3_X1 U17267 ( .A1(n26026), .A2(n26025), .A3(n23015), .ZN(n24030) );
  NOR3_X1 U17268 ( .A1(n26172), .A2(n24300), .A3(n24321), .ZN(n23018) );
  NOR2_X1 U17269 ( .A1(n26061), .A2(n24322), .ZN(n23020) );
  NAND3_X1 U17270 ( .A1(n25421), .A2(n24536), .A3(n25466), .ZN(n23021) );
  AND3_X1 U17271 ( .A1(n23020), .A2(n23019), .A3(n23018), .ZN(n23017) );
  MUX2_X1 U17272 ( .A(net713892), .B(n26136), .S(n24204), .Z(n23016) );
  NOR2_X1 U17273 ( .A1(n26135), .A2(net749977), .ZN(net714413) );
  OAI22_X1 U17274 ( .A1(n25448), .A2(net713897), .B1(n24030), .B2(net713882), 
        .ZN(net714414) );
  MUX2_X1 U17275 ( .A(net713728), .B(net717087), .S(n24204), .Z(net714410) );
  NOR2_X1 U17276 ( .A1(net749894), .A2(n23016), .ZN(net714409) );
  OAI22_X1 U17277 ( .A1(net742259), .A2(net750287), .B1(n24560), .B2(net718355), .ZN(net714434) );
  OAI222_X1 U17278 ( .A1(net717075), .A2(net749454), .B1(net728314), .B2(
        net718391), .C1(n24270), .C2(net713810), .ZN(net714432) );
  OAI222_X1 U17279 ( .A1(net717055), .A2(net742508), .B1(net762753), .B2(
        n25586), .C1(n25443), .C2(net713773), .ZN(net714433) );
  CLKBUF_X1 U17280 ( .A(net728481), .Z(net780602) );
  NAND2_X1 U17281 ( .A1(n22873), .A2(net787518), .ZN(net780598) );
  INV_X1 U17282 ( .A(n24357), .ZN(n23022) );
  CLKBUF_X3 U17283 ( .A(n25663), .Z(n24357) );
  AND2_X1 U17284 ( .A1(net749830), .A2(n23024), .ZN(n23909) );
  NOR3_X1 U17285 ( .A1(n23906), .A2(n26119), .A3(net714547), .ZN(n23024) );
  NOR2_X1 U17286 ( .A1(net741959), .A2(n4406), .ZN(n23025) );
  INV_X1 U17287 ( .A(net742017), .ZN(net780584) );
  OR2_X1 U17288 ( .A1(net717543), .A2(n24400), .ZN(n24291) );
  AND2_X2 U17289 ( .A1(net755056), .A2(net755048), .ZN(n24550) );
  NOR2_X1 U17290 ( .A1(net767335), .A2(n23933), .ZN(net780578) );
  BUF_X1 U17291 ( .A(net736739), .Z(net780579) );
  NOR3_X1 U17292 ( .A1(n23771), .A2(net342960), .A3(net342852), .ZN(net736739)
         );
  CLKBUF_X1 U17293 ( .A(net714873), .Z(net755075) );
  CLKBUF_X1 U17294 ( .A(n26110), .Z(n23027) );
  CLKBUF_X1 U17295 ( .A(net715176), .Z(net780568) );
  BUF_X1 U17296 ( .A(net718152), .Z(net742241) );
  CLKBUF_X1 U17297 ( .A(net718152), .Z(net749697) );
  NAND2_X1 U17298 ( .A1(net765341), .A2(n22684), .ZN(n26602) );
  NAND2_X1 U17299 ( .A1(n22851), .A2(n24395), .ZN(n23028) );
  BUF_X1 U17300 ( .A(net750277), .Z(net780556) );
  NOR2_X1 U17301 ( .A1(net715359), .A2(n23865), .ZN(n23029) );
  CLKBUF_X1 U17302 ( .A(net713753), .Z(net749812) );
  AOI221_X4 U17303 ( .B1(n25790), .B2(net732762), .C1(n23242), .C2(net732762), 
        .A(net780551), .ZN(n23243) );
  INV_X1 U17304 ( .A(net755238), .ZN(net780543) );
  OR2_X1 U17305 ( .A1(n24403), .A2(n24317), .ZN(n24339) );
  CLKBUF_X1 U17306 ( .A(n25415), .Z(n23030) );
  CLKBUF_X1 U17307 ( .A(net734282), .Z(net780528) );
  NAND3_X1 U17308 ( .A1(net714476), .A2(n24300), .A3(n24206), .ZN(n25774) );
  AND2_X1 U17309 ( .A1(n26269), .A2(n26268), .ZN(n23031) );
  NOR2_X1 U17310 ( .A1(n23031), .A2(net716311), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_5/N3 ) );
  OR2_X1 U17311 ( .A1(n19264), .A2(n19244), .ZN(n18346) );
  AND2_X1 U17312 ( .A1(n23779), .A2(n23780), .ZN(net712494) );
  INV_X1 U17313 ( .A(n25449), .ZN(n23295) );
  AND4_X1 U17314 ( .A1(n23282), .A2(n24611), .A3(n24583), .A4(n24581), .ZN(
        n26777) );
  BUF_X2 U17315 ( .A(net713866), .Z(net717056) );
  AND3_X1 U17316 ( .A1(net732754), .A2(n25413), .A3(n23368), .ZN(n25316) );
  OR2_X1 U17317 ( .A1(n23993), .A2(n1690), .ZN(n25506) );
  BUF_X1 U17318 ( .A(n26165), .Z(n25577) );
  INV_X1 U17319 ( .A(n25997), .ZN(n23713) );
  INV_X1 U17320 ( .A(n25922), .ZN(n25924) );
  OAI22_X1 U17321 ( .A1(n19395), .A2(n2926), .B1(n19383), .B2(n2929), .ZN(
        n23041) );
  OAI22_X1 U17322 ( .A1(n19385), .A2(n2925), .B1(n25267), .B2(n26785), .ZN(
        n23042) );
  AOI211_X1 U17323 ( .C1(n19530), .C2(n24690), .A(n23041), .B(n23042), .ZN(
        n23043) );
  AOI22_X1 U17324 ( .A1(n19337), .A2(n17831), .B1(n19336), .B2(n24709), .ZN(
        n23044) );
  AOI22_X1 U17325 ( .A1(n19373), .A2(n17836), .B1(n19372), .B2(n17837), .ZN(
        n23045) );
  NAND3_X1 U17326 ( .A1(n23043), .A2(n23044), .A3(n23045), .ZN(n25546) );
  AOI22_X1 U17327 ( .A1(n18347), .A2(n457), .B1(n451), .B2(net716461), .ZN(
        n23046) );
  OAI21_X1 U17328 ( .B1(net767169), .B2(n462), .A(n23046), .ZN(n23047) );
  AOI22_X1 U17329 ( .A1(n24767), .A2(net741532), .B1(n454), .B2(net741539), 
        .ZN(n23048) );
  OAI21_X1 U17330 ( .B1(n18332), .B2(n468), .A(n23048), .ZN(n23049) );
  AOI22_X1 U17331 ( .A1(n452), .A2(n18339), .B1(n455), .B2(n18338), .ZN(n23050) );
  AOI22_X1 U17332 ( .A1(net716491), .A2(n24766), .B1(n446), .B2(n18343), .ZN(
        n23051) );
  NAND2_X1 U17333 ( .A1(n23050), .A2(n23051), .ZN(n23052) );
  AOI22_X1 U17334 ( .A1(n18331), .A2(n17698), .B1(n453), .B2(n18330), .ZN(
        n23053) );
  AOI22_X1 U17335 ( .A1(n24769), .A2(net716417), .B1(n448), .B2(net767167), 
        .ZN(n23054) );
  AOI22_X1 U17336 ( .A1(n24768), .A2(net767214), .B1(n17697), .B2(n18328), 
        .ZN(n23055) );
  OAI22_X1 U17337 ( .A1(n18394), .A2(n24656), .B1(n463), .B2(net741541), .ZN(
        n23056) );
  OAI22_X1 U17338 ( .A1(n18395), .A2(n24655), .B1(n474), .B2(net741544), .ZN(
        n23057) );
  OAI22_X1 U17339 ( .A1(n18388), .A2(n475), .B1(n1755), .B2(net741549), .ZN(
        n23058) );
  OAI22_X1 U17340 ( .A1(n18318), .A2(n24654), .B1(n465), .B2(net518461), .ZN(
        n23059) );
  OAI22_X1 U17341 ( .A1(n18316), .A2(n472), .B1(n18315), .B2(n473), .ZN(n23060) );
  AOI211_X1 U17342 ( .C1(n18312), .C2(n459), .A(n23059), .B(n23060), .ZN(
        n23061) );
  AOI22_X1 U17343 ( .A1(n18310), .A2(n461), .B1(n18311), .B2(n447), .ZN(n23062) );
  AOI22_X1 U17344 ( .A1(n18321), .A2(n458), .B1(n456), .B2(net767173), .ZN(
        n23063) );
  NAND3_X1 U17345 ( .A1(n23061), .A2(n23062), .A3(n23063), .ZN(n23064) );
  NOR4_X1 U17346 ( .A1(n23056), .A2(n23057), .A3(n23058), .A4(n23064), .ZN(
        n23065) );
  NAND4_X1 U17347 ( .A1(n23053), .A2(n23054), .A3(n23055), .A4(n23065), .ZN(
        n23066) );
  NOR4_X1 U17348 ( .A1(n23047), .A2(n23049), .A3(n23052), .A4(n23066), .ZN(
        n23067) );
  NAND3_X1 U17349 ( .A1(n19644), .A2(n19642), .A3(n19643), .ZN(n23068) );
  NAND3_X1 U17350 ( .A1(n19647), .A2(n19646), .A3(n19641), .ZN(n23069) );
  NOR4_X1 U17351 ( .A1(n26332), .A2(n26331), .A3(n23068), .A4(n23069), .ZN(
        n23070) );
  NOR2_X1 U17352 ( .A1(n26637), .A2(n23070), .ZN(n23071) );
  OAI221_X1 U17353 ( .B1(n23071), .B2(n25665), .C1(n23071), .C2(n26603), .A(
        net716243), .ZN(n26333) );
  OAI22_X1 U17354 ( .A1(n19395), .A2(n2998), .B1(n3001), .B2(n19383), .ZN(
        n23072) );
  OAI22_X1 U17355 ( .A1(n19385), .A2(n2997), .B1(n24842), .B2(n26785), .ZN(
        n23073) );
  AOI211_X1 U17356 ( .C1(n19530), .C2(n24681), .A(n23072), .B(n23073), .ZN(
        n23074) );
  AOI22_X1 U17357 ( .A1(n19373), .A2(n17853), .B1(n19372), .B2(n17854), .ZN(
        n23075) );
  AOI22_X1 U17358 ( .A1(n19337), .A2(n17848), .B1(n19336), .B2(n24682), .ZN(
        n23076) );
  NAND3_X1 U17359 ( .A1(n23074), .A2(n23075), .A3(n23076), .ZN(n26666) );
  OAI22_X1 U17360 ( .A1(net716477), .A2(n2304), .B1(net767232), .B2(n24623), 
        .ZN(n23077) );
  OAI22_X1 U17361 ( .A1(n18362), .A2(n2300), .B1(n18361), .B2(n2301), .ZN(
        n23078) );
  OAI22_X1 U17362 ( .A1(n24594), .A2(n18332), .B1(net767172), .B2(n2306), .ZN(
        n23079) );
  OAI22_X1 U17363 ( .A1(n18401), .A2(n2297), .B1(n18400), .B2(n2314), .ZN(
        n23080) );
  OAI22_X1 U17364 ( .A1(net767237), .A2(n24675), .B1(n18369), .B2(n2303), .ZN(
        n23081) );
  NOR2_X1 U17365 ( .A1(n23080), .A2(n23081), .ZN(n23082) );
  OAI21_X1 U17366 ( .B1(n24676), .B2(n18363), .A(n23082), .ZN(n23083) );
  NOR4_X1 U17367 ( .A1(n23077), .A2(n23078), .A3(n23079), .A4(n23083), .ZN(
        n23084) );
  OAI22_X1 U17368 ( .A1(n18393), .A2(n2319), .B1(n18394), .B2(n2316), .ZN(
        n23085) );
  AOI22_X1 U17369 ( .A1(n18001), .A2(net767235), .B1(n17991), .B2(net716417), 
        .ZN(n23086) );
  OAI22_X1 U17370 ( .A1(n18318), .A2(n2298), .B1(n18390), .B2(n2313), .ZN(
        n23087) );
  OAI22_X1 U17371 ( .A1(n18388), .A2(n24674), .B1(n18387), .B2(n2317), .ZN(
        n23088) );
  AOI211_X1 U17372 ( .C1(net716405), .C2(n18000), .A(n23087), .B(n23088), .ZN(
        n23089) );
  OAI211_X1 U17373 ( .C1(n18395), .C2(n2322), .A(n23086), .B(n23089), .ZN(
        n23090) );
  AOI211_X1 U17374 ( .C1(n17990), .C2(net767239), .A(n23085), .B(n23090), .ZN(
        n23091) );
  OAI211_X1 U17375 ( .C1(n18382), .C2(n2320), .A(n23084), .B(n23091), .ZN(
        n25527) );
  NAND3_X1 U17376 ( .A1(n19842), .A2(n19840), .A3(n19841), .ZN(n23092) );
  NOR4_X1 U17377 ( .A1(n26636), .A2(n26635), .A3(n26634), .A4(n23092), .ZN(
        n23093) );
  NOR2_X1 U17378 ( .A1(n26637), .A2(n23093), .ZN(n23094) );
  OAI221_X1 U17379 ( .B1(n23094), .B2(net717048), .C1(n23094), .C2(n26706), 
        .A(net716243), .ZN(n26638) );
  NAND2_X1 U17380 ( .A1(n20084), .A2(n20061), .ZN(n19350) );
  NAND2_X1 U17381 ( .A1(n25502), .A2(net749289), .ZN(n23095) );
  OAI21_X1 U17382 ( .B1(n23096), .B2(n26563), .A(n26565), .ZN(n23097) );
  OAI21_X1 U17383 ( .B1(n23097), .B2(n25366), .A(n26566), .ZN(n23098) );
  NAND2_X1 U17384 ( .A1(n23098), .A2(net717091), .ZN(n23099) );
  AOI21_X1 U17385 ( .B1(n24529), .B2(n23095), .A(net712880), .ZN(n23100) );
  OAI21_X1 U17386 ( .B1(n23023), .B2(n23100), .A(n26560), .ZN(n23101) );
  NAND2_X1 U17387 ( .A1(net755683), .A2(net755757), .ZN(n23102) );
  OAI21_X1 U17388 ( .B1(net712855), .B2(n23102), .A(net732762), .ZN(n23103) );
  OAI221_X1 U17389 ( .B1(n23099), .B2(n26562), .C1(n23099), .C2(n23101), .A(
        n23103), .ZN(n23104) );
  AOI22_X1 U17390 ( .A1(n726), .A2(n19336), .B1(n24800), .B2(n19393), .ZN(
        n23105) );
  OAI21_X1 U17391 ( .B1(n741), .B2(n19338), .A(n23105), .ZN(n23106) );
  AOI22_X1 U17392 ( .A1(n733), .A2(n19314), .B1(n24692), .B2(n23994), .ZN(
        n23107) );
  AOI22_X1 U17393 ( .A1(n17748), .A2(n25683), .B1(n17749), .B2(n19315), .ZN(
        n23108) );
  AOI22_X1 U17394 ( .A1(n720), .A2(n19319), .B1(n734), .B2(n19318), .ZN(n23109) );
  OAI22_X1 U17395 ( .A1(n745), .A2(n19324), .B1(n746), .B2(n19323), .ZN(n23110) );
  AOI22_X1 U17396 ( .A1(n19327), .A2(n729), .B1(n731), .B2(n19328), .ZN(n23111) );
  AOI22_X1 U17397 ( .A1(n723), .A2(n19530), .B1(n732), .B2(n19320), .ZN(n23112) );
  OAI211_X1 U17398 ( .C1(n738), .C2(n26785), .A(n23111), .B(n23112), .ZN(
        n23113) );
  AOI22_X1 U17399 ( .A1(n725), .A2(n19345), .B1(n728), .B2(n19344), .ZN(n23114) );
  NOR2_X1 U17400 ( .A1(n25678), .A2(n24624), .ZN(n23115) );
  OAI22_X1 U17401 ( .A1(n743), .A2(n25675), .B1(n744), .B2(n25677), .ZN(n23116) );
  AOI211_X1 U17402 ( .C1(n19348), .C2(n719), .A(n23115), .B(n23116), .ZN(
        n23117) );
  AOI22_X1 U17403 ( .A1(n730), .A2(n19351), .B1(n724), .B2(n25679), .ZN(n23118) );
  NAND3_X1 U17404 ( .A1(n23114), .A2(n23117), .A3(n23118), .ZN(n23119) );
  AOI22_X1 U17405 ( .A1(n24742), .A2(n23995), .B1(n722), .B2(n19308), .ZN(
        n23120) );
  AOI22_X1 U17406 ( .A1(n24741), .A2(n19333), .B1(n721), .B2(n24026), .ZN(
        n23121) );
  AOI22_X1 U17407 ( .A1(n17747), .A2(n25681), .B1(n17745), .B2(n24007), .ZN(
        n23122) );
  NAND3_X1 U17408 ( .A1(n23120), .A2(n23121), .A3(n23122), .ZN(n23123) );
  NOR4_X1 U17409 ( .A1(n23110), .A2(n23113), .A3(n23119), .A4(n23123), .ZN(
        n23124) );
  NAND4_X1 U17410 ( .A1(n23107), .A2(n23108), .A3(n23109), .A4(n23124), .ZN(
        n23125) );
  AOI211_X1 U17411 ( .C1(n17746), .C2(n19337), .A(n23106), .B(n23125), .ZN(
        n26456) );
  NAND4_X1 U17412 ( .A1(n18335), .A2(n18337), .A3(n18336), .A4(n26681), .ZN(
        n23126) );
  NOR3_X1 U17413 ( .A1(n26683), .A2(n23126), .A3(n26682), .ZN(n23127) );
  NOR2_X1 U17414 ( .A1(n23127), .A2(n24008), .ZN(n23128) );
  OAI221_X1 U17415 ( .B1(n23128), .B2(net712397), .C1(n23128), .C2(n26684), 
        .A(net742649), .ZN(n26685) );
  AOI222_X1 U17416 ( .A1(n18372), .A2(n17935), .B1(n14127), .B2(net712520), 
        .C1(n17928), .C2(net716423), .ZN(n23129) );
  AOI222_X1 U17417 ( .A1(net767238), .A2(n17925), .B1(n24738), .B2(net716461), 
        .C1(n24597), .C2(net767167), .ZN(n23130) );
  AOI22_X1 U17418 ( .A1(n18373), .A2(n17934), .B1(net767214), .B2(n17931), 
        .ZN(n23131) );
  AND3_X1 U17419 ( .A1(n23129), .A2(n23130), .A3(n23131), .ZN(n24046) );
  OAI211_X1 U17420 ( .C1(n468), .C2(n19338), .A(n26359), .B(n19511), .ZN(
        n23132) );
  NAND3_X1 U17421 ( .A1(n19514), .A2(n19512), .A3(n19513), .ZN(n23133) );
  NOR4_X1 U17422 ( .A1(n26361), .A2(n26360), .A3(n23132), .A4(n23133), .ZN(
        n23134) );
  NOR2_X1 U17423 ( .A1(n26637), .A2(n23134), .ZN(n23135) );
  OAI221_X1 U17424 ( .B1(n23135), .B2(net712499), .C1(n23135), .C2(n26662), 
        .A(net716259), .ZN(n26362) );
  NAND3_X1 U17425 ( .A1(net717074), .A2(net728314), .A3(net712469), .ZN(n23136) );
  NOR4_X1 U17426 ( .A1(net712467), .A2(net712468), .A3(net712466), .A4(n23136), 
        .ZN(n23137) );
  AOI21_X1 U17427 ( .B1(net712462), .B2(n23137), .A(net729186), .ZN(n23138) );
  OAI21_X1 U17428 ( .B1(net713154), .B2(net741975), .A(net712472), .ZN(n23139)
         );
  NAND3_X1 U17429 ( .A1(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [20]), .A2(net712795), .A3(net780360), .ZN(net712812) );
  NOR2_X1 U17430 ( .A1(n18394), .A2(n2928), .ZN(n23140) );
  OAI22_X1 U17431 ( .A1(n18382), .A2(n2932), .B1(n18393), .B2(n2931), .ZN(
        n23141) );
  AOI211_X1 U17432 ( .C1(net767239), .C2(n17827), .A(n23140), .B(n23141), .ZN(
        n23142) );
  AOI22_X1 U17433 ( .A1(n18307), .A2(n17840), .B1(n17838), .B2(net716405), 
        .ZN(n23143) );
  AOI22_X1 U17434 ( .A1(n17833), .A2(net767214), .B1(n17830), .B2(net716423), 
        .ZN(n23144) );
  OAI22_X1 U17435 ( .A1(net767172), .A2(n2918), .B1(n2919), .B2(n18346), .ZN(
        n23145) );
  OAI22_X1 U17436 ( .A1(n18367), .A2(n24637), .B1(n2909), .B2(n18401), .ZN(
        n23146) );
  OAI22_X1 U17437 ( .A1(net767237), .A2(n24638), .B1(n2916), .B2(net716477), 
        .ZN(n23147) );
  OAI22_X1 U17438 ( .A1(n18369), .A2(n2915), .B1(n2913), .B2(n18361), .ZN(
        n23148) );
  NOR4_X1 U17439 ( .A1(n23145), .A2(n23146), .A3(n23147), .A4(n23148), .ZN(
        n23149) );
  AOI22_X1 U17440 ( .A1(n17839), .A2(net767235), .B1(n24711), .B2(n18300), 
        .ZN(n23150) );
  AOI22_X1 U17441 ( .A1(n17828), .A2(n18326), .B1(n24710), .B2(net767167), 
        .ZN(n23151) );
  AOI22_X1 U17442 ( .A1(net767238), .A2(n17826), .B1(n17832), .B2(net767171), 
        .ZN(n23152) );
  AND4_X1 U17443 ( .A1(n23149), .A2(n23150), .A3(n23151), .A4(n23152), .ZN(
        n23153) );
  AND4_X1 U17444 ( .A1(n23142), .A2(n23143), .A3(n23144), .A4(n23153), .ZN(
        n26701) );
  OAI211_X1 U17445 ( .C1(n19338), .C2(n976), .A(n26325), .B(n19887), .ZN(
        n23154) );
  NAND3_X1 U17446 ( .A1(n19886), .A2(n19884), .A3(n19885), .ZN(n23155) );
  NAND3_X1 U17447 ( .A1(n19889), .A2(n19888), .A3(n19883), .ZN(n23156) );
  NOR4_X1 U17448 ( .A1(n26326), .A2(n23154), .A3(n23155), .A4(n23156), .ZN(
        n23157) );
  NOR2_X1 U17449 ( .A1(n26637), .A2(n23157), .ZN(n23158) );
  OAI221_X1 U17450 ( .B1(n23158), .B2(net712499), .C1(n23158), .C2(n26327), 
        .A(net716255), .ZN(n26328) );
  NAND2_X1 U17451 ( .A1(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [26]), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [27]), .ZN(net780340) );
  INV_X1 U17452 ( .A(net732762), .ZN(net780337) );
  AOI22_X1 U17453 ( .A1(n339), .A2(n25679), .B1(n24801), .B2(n19393), .ZN(
        n23159) );
  OAI21_X1 U17454 ( .B1(n356), .B2(n19338), .A(n23159), .ZN(n23160) );
  AOI22_X1 U17455 ( .A1(n17679), .A2(n19335), .B1(n17677), .B2(n19334), .ZN(
        n23161) );
  AOI22_X1 U17456 ( .A1(n24772), .A2(n25682), .B1(n336), .B2(n24026), .ZN(
        n23162) );
  AOI22_X1 U17457 ( .A1(n17678), .A2(n19337), .B1(n341), .B2(n19336), .ZN(
        n23163) );
  AOI22_X1 U17458 ( .A1(n17680), .A2(n25683), .B1(n17681), .B2(n19315), .ZN(
        n23164) );
  OAI21_X1 U17459 ( .B1(n351), .B2(n24614), .A(n23164), .ZN(n23165) );
  AOI22_X1 U17460 ( .A1(n348), .A2(n19314), .B1(n19308), .B2(n337), .ZN(n23166) );
  OAI21_X1 U17461 ( .B1(n363), .B2(n24613), .A(n23166), .ZN(n23167) );
  AOI22_X1 U17462 ( .A1(n19327), .A2(n344), .B1(n19328), .B2(n346), .ZN(n23168) );
  AOI22_X1 U17463 ( .A1(n335), .A2(n19319), .B1(n349), .B2(n19318), .ZN(n23169) );
  OAI22_X1 U17464 ( .A1(n19326), .A2(n24667), .B1(n353), .B2(n26785), .ZN(
        n23170) );
  OAI22_X1 U17465 ( .A1(n19324), .A2(n360), .B1(n361), .B2(n19323), .ZN(n23171) );
  AOI211_X1 U17466 ( .C1(n19320), .C2(n347), .A(n23170), .B(n23171), .ZN(
        n23172) );
  NAND3_X1 U17467 ( .A1(n23168), .A2(n23169), .A3(n23172), .ZN(n23173) );
  AOI22_X1 U17468 ( .A1(n24771), .A2(n24591), .B1(n342), .B2(n24617), .ZN(
        n23174) );
  AOI22_X1 U17469 ( .A1(n340), .A2(n19345), .B1(n343), .B2(n19344), .ZN(n23175) );
  AOI22_X1 U17470 ( .A1(n24770), .A2(n24619), .B1(n334), .B2(n19348), .ZN(
        n23176) );
  NAND3_X1 U17471 ( .A1(n23174), .A2(n23175), .A3(n23176), .ZN(n23177) );
  NOR4_X1 U17472 ( .A1(n23165), .A2(n23167), .A3(n23173), .A4(n23177), .ZN(
        n23178) );
  NAND4_X1 U17473 ( .A1(n23161), .A2(n23162), .A3(n23163), .A4(n23178), .ZN(
        n23179) );
  AOI211_X1 U17474 ( .C1(n345), .C2(n25667), .A(n23160), .B(n23179), .ZN(
        n26505) );
  AOI22_X1 U17475 ( .A1(n18310), .A2(n929), .B1(n18311), .B2(n915), .ZN(n23180) );
  AOI22_X1 U17476 ( .A1(n18306), .A2(n928), .B1(net767239), .B2(n24691), .ZN(
        n23181) );
  AOI22_X1 U17477 ( .A1(n18307), .A2(n17783), .B1(net716405), .B2(n17782), 
        .ZN(n23182) );
  AOI22_X1 U17478 ( .A1(n18347), .A2(n925), .B1(net716461), .B2(n919), .ZN(
        n23183) );
  NAND4_X1 U17479 ( .A1(n23180), .A2(n23181), .A3(n23182), .A4(n23183), .ZN(
        n23184) );
  OAI22_X1 U17480 ( .A1(n18316), .A2(n940), .B1(n18315), .B2(n941), .ZN(n23185) );
  AOI22_X1 U17481 ( .A1(n18321), .A2(n926), .B1(net767173), .B2(n924), .ZN(
        n23186) );
  AOI22_X1 U17482 ( .A1(n18529), .A2(n918), .B1(n18312), .B2(n927), .ZN(n23187) );
  OAI211_X1 U17483 ( .C1(n933), .C2(net518461), .A(n23186), .B(n23187), .ZN(
        n23188) );
  AOI22_X1 U17484 ( .A1(n18339), .A2(n920), .B1(n18338), .B2(n923), .ZN(n23189) );
  OAI22_X1 U17485 ( .A1(net767237), .A2(n938), .B1(n939), .B2(net767232), .ZN(
        n23190) );
  AOI21_X1 U17486 ( .B1(n914), .B2(n18343), .A(n23190), .ZN(n23191) );
  OAI211_X1 U17487 ( .C1(net716477), .C2(n24622), .A(n23189), .B(n23191), .ZN(
        n23192) );
  OR4_X1 U17488 ( .A1(n23184), .A2(n23185), .A3(n23188), .A4(n23192), .ZN(
        n25571) );
  NAND3_X1 U17489 ( .A1(net716247), .A2(n25335), .A3(n18136), .ZN(n23194) );
  NAND3_X1 U17490 ( .A1(n23193), .A2(n23194), .A3(n22742), .ZN(
        \core_inst/IDEX_RF_ADDR_DEST/DFF_0/N3 ) );
  NOR2_X1 U17491 ( .A1(n5577), .A2(n24343), .ZN(n23195) );
  NAND3_X1 U17492 ( .A1(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [10]), .A2(n26575), .A3(n23195), .ZN(n26573) );
  INV_X1 U17493 ( .A(net712795), .ZN(net780298) );
  INV_X1 U17494 ( .A(net780602), .ZN(net780291) );
  NAND3_X1 U17495 ( .A1(net749442), .A2(n26256), .A3(net749719), .ZN(n23196)
         );
  OAI211_X1 U17496 ( .C1(n24530), .C2(n23196), .A(net713463), .B(net755052), 
        .ZN(net780293) );
  AOI22_X1 U17497 ( .A1(n842), .A2(n19345), .B1(n845), .B2(n19344), .ZN(n23197) );
  AOI22_X1 U17498 ( .A1(n847), .A2(n19351), .B1(n841), .B2(n25679), .ZN(n23198) );
  NAND2_X1 U17499 ( .A1(n836), .A2(n19348), .ZN(n23199) );
  OAI21_X1 U17500 ( .B1(n861), .B2(n25677), .A(n23199), .ZN(n23200) );
  OAI22_X1 U17501 ( .A1(n25678), .A2(net741520), .B1(n860), .B2(n25675), .ZN(
        n23201) );
  OAI22_X1 U17502 ( .A1(n862), .A2(n19324), .B1(n863), .B2(n19323), .ZN(n23202) );
  AOI22_X1 U17503 ( .A1(n19327), .A2(n846), .B1(n848), .B2(n19328), .ZN(n23203) );
  AOI22_X1 U17504 ( .A1(n840), .A2(n19530), .B1(n849), .B2(n19320), .ZN(n23204) );
  OAI211_X1 U17505 ( .C1(n855), .C2(n26785), .A(n23203), .B(n23204), .ZN(
        n23205) );
  NOR4_X1 U17506 ( .A1(n23200), .A2(n23201), .A3(n23202), .A4(n23205), .ZN(
        n23206) );
  NAND3_X1 U17507 ( .A1(n23197), .A2(n23198), .A3(n23206), .ZN(n26516) );
  NAND2_X1 U17508 ( .A1(n26405), .A2(n24830), .ZN(n23207) );
  NAND3_X1 U17509 ( .A1(n26404), .A2(net713168), .A3(net740526), .ZN(n23208)
         );
  AOI21_X1 U17510 ( .B1(net749830), .B2(n23208), .A(net713167), .ZN(n23209) );
  OAI21_X1 U17511 ( .B1(n24297), .B2(n23209), .A(net755714), .ZN(n23210) );
  XNOR2_X1 U17512 ( .A(n23210), .B(n23207), .ZN(n23211) );
  OAI211_X1 U17513 ( .C1(net713154), .C2(n23211), .A(n26407), .B(n26406), .ZN(
        n23212) );
  INV_X1 U17514 ( .A(n26408), .ZN(n23213) );
  INV_X1 U17515 ( .A(net749936), .ZN(net780262) );
  OAI221_X1 U17516 ( .B1(net749936), .B2(n23213), .C1(net780262), .C2(
        net713152), .A(net713148), .ZN(n23214) );
  NOR3_X1 U17517 ( .A1(n23305), .A2(n23212), .A3(n23214), .ZN(n26735) );
  NAND3_X1 U17518 ( .A1(net755708), .A2(net718074), .A3(s_IFID_IR[18]), .ZN(
        n23215) );
  NAND3_X1 U17519 ( .A1(n23215), .A2(n22742), .A3(n23216), .ZN(
        \core_inst/IDEX_RF_ADDR_DEST/DFF_2/N3 ) );
  NOR3_X1 U17520 ( .A1(n25933), .A2(n25338), .A3(net713442), .ZN(n26732) );
  AOI22_X1 U17521 ( .A1(n19315), .A2(n17891), .B1(n17889), .B2(n25683), .ZN(
        n23217) );
  NOR2_X1 U17522 ( .A1(n3075), .A2(n19388), .ZN(n23218) );
  OAI22_X1 U17523 ( .A1(n19389), .A2(n3072), .B1(n19378), .B2(n3076), .ZN(
        n23219) );
  AOI211_X1 U17524 ( .C1(n17878), .C2(n23994), .A(n23218), .B(n23219), .ZN(
        n23220) );
  AOI22_X1 U17525 ( .A1(n17890), .A2(n23995), .B1(n24703), .B2(n19308), .ZN(
        n23221) );
  OAI22_X1 U17526 ( .A1(n3062), .A2(n26614), .B1(n3063), .B2(n19350), .ZN(
        n23222) );
  OAI22_X1 U17527 ( .A1(n25677), .A2(n24631), .B1(n3053), .B2(n19396), .ZN(
        n23223) );
  OAI22_X1 U17528 ( .A1(n25678), .A2(n3060), .B1(n25676), .B2(n24632), .ZN(
        n23224) );
  OAI22_X1 U17529 ( .A1(n19365), .A2(n3057), .B1(n19370), .B2(n3059), .ZN(
        n23225) );
  NOR4_X1 U17530 ( .A1(n23222), .A2(n23223), .A3(n23224), .A4(n23225), .ZN(
        n23226) );
  NAND4_X1 U17531 ( .A1(n23217), .A2(n23220), .A3(n23221), .A4(n23226), .ZN(
        n26629) );
  AOI22_X1 U17532 ( .A1(net716417), .A2(n17960), .B1(n24727), .B2(net767167), 
        .ZN(n23227) );
  AOI22_X1 U17533 ( .A1(net767238), .A2(n17958), .B1(n14393), .B2(net767171), 
        .ZN(n23228) );
  AOI22_X1 U17534 ( .A1(net767214), .A2(n17963), .B1(n17961), .B2(n18328), 
        .ZN(n23229) );
  OAI22_X1 U17535 ( .A1(net767172), .A2(n2162), .B1(n2163), .B2(n18346), .ZN(
        n23230) );
  OAI22_X1 U17536 ( .A1(net767232), .A2(n24775), .B1(n2153), .B2(n18401), .ZN(
        n23231) );
  OAI22_X1 U17537 ( .A1(net716477), .A2(n2160), .B1(net767237), .B2(n24776), 
        .ZN(n23232) );
  OAI22_X1 U17538 ( .A1(n18361), .A2(n2157), .B1(n18369), .B2(n2159), .ZN(
        n23233) );
  NOR4_X1 U17539 ( .A1(n23230), .A2(n23231), .A3(n23232), .A4(n23233), .ZN(
        n23234) );
  AND4_X1 U17540 ( .A1(n23227), .A2(n23228), .A3(n23229), .A4(n23234), .ZN(
        n23235) );
  AOI22_X1 U17541 ( .A1(n18307), .A2(n17970), .B1(n17968), .B2(net716405), 
        .ZN(n23236) );
  NOR2_X1 U17542 ( .A1(n18393), .A2(n2175), .ZN(n23237) );
  OAI22_X1 U17543 ( .A1(n18382), .A2(n2176), .B1(n18394), .B2(n2172), .ZN(
        n23238) );
  AOI211_X1 U17544 ( .C1(net767239), .C2(n17959), .A(n23237), .B(n23238), .ZN(
        n23239) );
  AOI22_X1 U17545 ( .A1(n18300), .A2(n24728), .B1(n17969), .B2(net767235), 
        .ZN(n23240) );
  NAND4_X1 U17546 ( .A1(n23235), .A2(n23236), .A3(n23239), .A4(n23240), .ZN(
        n25567) );
  NAND3_X1 U17547 ( .A1(n14191), .A2(s_IFID_IR[27]), .A3(n24611), .ZN(n23241)
         );
  OR3_X1 U17548 ( .A1(s_IFID_IR[29]), .A2(n18138), .A3(n23241), .ZN(n18133) );
  XOR2_X1 U17549 ( .A(net712847), .B(n6180), .Z(n26568) );
  INV_X1 U17550 ( .A(n26120), .ZN(n23242) );
  NAND2_X1 U17551 ( .A1(net796204), .A2(n23243), .ZN(n23298) );
  AOI21_X1 U17552 ( .B1(n26428), .B2(n25665), .A(n26429), .ZN(n23244) );
  NOR2_X1 U17553 ( .A1(n23244), .A2(net785239), .ZN(
        \core_inst/IDEX_RF_IN1/DFF_19/N3 ) );
  NAND2_X1 U17554 ( .A1(n24398), .A2(n24397), .ZN(n23245) );
  NOR3_X1 U17555 ( .A1(n24399), .A2(n24234), .A3(n23245), .ZN(n24334) );
  NAND2_X1 U17556 ( .A1(net758544), .A2(net714239), .ZN(n23246) );
  NOR2_X1 U17557 ( .A1(n23290), .A2(n23246), .ZN(n26728) );
  AOI222_X1 U17558 ( .A1(net740710), .A2(net741608), .B1(net712606), .B2(
        n24811), .C1(n17858), .C2(n26663), .ZN(n23247) );
  INV_X1 U17559 ( .A(n23247), .ZN(n26714) );
  NOR2_X1 U17560 ( .A1(net738518), .A2(net780214), .ZN(n26738) );
  OAI22_X1 U17561 ( .A1(n19395), .A2(n3070), .B1(n19383), .B2(n3073), .ZN(
        n23248) );
  OAI22_X1 U17562 ( .A1(n19385), .A2(n3069), .B1(n25265), .B2(n26785), .ZN(
        n23249) );
  AOI211_X1 U17563 ( .C1(n19530), .C2(n24688), .A(n23248), .B(n23249), .ZN(
        n23250) );
  AOI22_X1 U17564 ( .A1(n19337), .A2(n17882), .B1(n19336), .B2(n24701), .ZN(
        n23251) );
  AOI22_X1 U17565 ( .A1(n19373), .A2(n17887), .B1(n19372), .B2(n17888), .ZN(
        n23252) );
  NAND3_X1 U17566 ( .A1(n23250), .A2(n23251), .A3(n23252), .ZN(n26628) );
  OAI22_X1 U17567 ( .A1(n18400), .A2(n2170), .B1(n18387), .B2(n2173), .ZN(
        n23253) );
  OAI22_X1 U17568 ( .A1(n18390), .A2(n2169), .B1(net518461), .B2(n25326), .ZN(
        n23254) );
  AOI211_X1 U17569 ( .C1(n18529), .C2(n24788), .A(n23253), .B(n23254), .ZN(
        n23255) );
  AOI22_X1 U17570 ( .A1(n18331), .A2(n17962), .B1(n18330), .B2(n24789), .ZN(
        n23256) );
  AOI22_X1 U17571 ( .A1(n18373), .A2(n17966), .B1(n18372), .B2(n17967), .ZN(
        n23257) );
  NAND3_X1 U17572 ( .A1(n23255), .A2(n23256), .A3(n23257), .ZN(n25568) );
  AOI21_X1 U17573 ( .B1(net717091), .B2(net780528), .A(net742518), .ZN(n26730)
         );
  NOR3_X1 U17574 ( .A1(net713850), .A2(net713849), .A3(net749607), .ZN(n26734)
         );
  NOR2_X1 U17575 ( .A1(n6180), .A2(net712847), .ZN(n23258) );
  XNOR2_X1 U17576 ( .A(n23258), .B(n6546), .ZN(n26410) );
  NOR3_X1 U17577 ( .A1(n18196), .A2(net720303), .A3(n18143), .ZN(n23259) );
  NAND2_X1 U17578 ( .A1(net713389), .A2(n23259), .ZN(\cu_inst/EX/DFF_1/N3 ) );
  CLKBUF_X3 U17579 ( .A(net741307), .Z(net716221) );
  CLKBUF_X3 U17580 ( .A(net741307), .Z(net716223) );
  NAND2_X2 U17581 ( .A1(n20076), .A2(n20064), .ZN(n19338) );
  INV_X2 U17582 ( .A(n19350), .ZN(n25679) );
  OAI21_X2 U17583 ( .B1(net714586), .B2(n25972), .A(n24172), .ZN(net713966) );
  BUF_X2 U17584 ( .A(net717104), .Z(net717106) );
  AND2_X1 U17585 ( .A1(net742286), .A2(n24351), .ZN(n23262) );
  INV_X1 U17586 ( .A(n23272), .ZN(n26605) );
  OAI21_X1 U17587 ( .B1(n26604), .B2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [4]), .A(n26710), .ZN(n23272) );
  OAI211_X1 U17588 ( .C1(n18153), .C2(net741565), .A(n18159), .B(n18186), .ZN(
        \cu_inst/EX/DFF_12/N3 ) );
  NAND3_X1 U17589 ( .A1(n14128), .A2(n26777), .A3(n18162), .ZN(n18186) );
  INV_X1 U17590 ( .A(n23273), .ZN(n24168) );
  OAI21_X1 U17591 ( .B1(n26709), .B2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [6]), .A(n26671), .ZN(n23273) );
  OAI221_X1 U17592 ( .B1(n18139), .B2(n18140), .C1(n18139), .C2(n18141), .A(
        n18142), .ZN(\cu_inst/EX/DFF_17/N3 ) );
  NOR2_X1 U17593 ( .A1(n18143), .A2(net720303), .ZN(n18142) );
  NOR2_X1 U17594 ( .A1(n18145), .A2(n18146), .ZN(n18141) );
  OAI211_X1 U17595 ( .C1(n18139), .C2(n18173), .A(n18164), .B(n18174), .ZN(
        \cu_inst/EX/DFF_13/N3 ) );
  OAI21_X1 U17596 ( .B1(n18175), .B2(n24813), .A(s_IFID_IR[30]), .ZN(n18174)
         );
  NAND4_X1 U17597 ( .A1(n18062), .A2(n14128), .A3(n18059), .A4(n24616), .ZN(
        n18173) );
  AOI211_X1 U17598 ( .C1(n18156), .C2(n18146), .A(n18177), .B(n18178), .ZN(
        n18164) );
  OAI211_X1 U17599 ( .C1(n18153), .C2(n18138), .A(n18179), .B(n18180), .ZN(
        n18178) );
  OAI221_X1 U17600 ( .B1(n18181), .B2(n18182), .C1(n18181), .C2(n14190), .A(
        n26777), .ZN(n18180) );
  NOR3_X1 U17601 ( .A1(n24584), .A2(net741565), .A3(n18171), .ZN(n18177) );
  NAND3_X1 U17602 ( .A1(net709330), .A2(n18148), .A3(n18129), .ZN(
        \cu_inst/EX/DFF_16/N3 ) );
  AOI211_X1 U17603 ( .C1(n26777), .C2(n18150), .A(n18151), .B(n18152), .ZN(
        n18148) );
  OAI21_X1 U17604 ( .B1(n23274), .B2(n26258), .A(net741565), .ZN(n18193) );
  NAND2_X1 U17605 ( .A1(n18129), .A2(n26779), .ZN(n23274) );
  NAND2_X1 U17606 ( .A1(n23275), .A2(n23276), .ZN(net713414) );
  NOR3_X1 U17607 ( .A1(n23277), .A2(n23278), .A3(n23279), .ZN(n23276) );
  NAND2_X1 U17608 ( .A1(s_ID_rf_write_en), .A2(n19290), .ZN(n23279) );
  AOI22_X1 U17609 ( .A1(s_IFID_IR[19]), .A2(n19288), .B1(s_IFID_IR[18]), .B2(
        n19289), .ZN(n19290) );
  INV_X1 U17610 ( .A(n19293), .ZN(n23278) );
  AOI22_X1 U17611 ( .A1(s_IFID_IR[20]), .A2(n19291), .B1(s_IFID_IR[17]), .B2(
        n19292), .ZN(n19293) );
  XNOR2_X1 U17612 ( .A(n19294), .B(s_IFID_IR[16]), .ZN(n23277) );
  NOR2_X1 U17613 ( .A1(n23280), .A2(n23281), .ZN(n23275) );
  OAI22_X1 U17614 ( .A1(s_IFID_IR[20]), .A2(n19291), .B1(n19288), .B2(
        s_IFID_IR[19]), .ZN(n23281) );
  OAI22_X1 U17615 ( .A1(s_IFID_IR[17]), .A2(n19292), .B1(n19289), .B2(
        s_IFID_IR[18]), .ZN(n23280) );
  INV_X1 U17616 ( .A(\core_inst/MEM/MUX_LOAD/MUX_BIT_12/s_top ), .ZN(n18223)
         );
  INV_X1 U17617 ( .A(\core_inst/MEM/MUX_LOAD/MUX_BIT_13/s_top ), .ZN(n18222)
         );
  INV_X1 U17618 ( .A(\core_inst/MEM/MUX_LOAD/MUX_BIT_14/s_top ), .ZN(n18221)
         );
  INV_X1 U17619 ( .A(\core_inst/MEM/MUX_LOAD/MUX_BIT_11/s_top ), .ZN(n18224)
         );
  INV_X1 U17620 ( .A(\core_inst/MEM/MUX_LOAD/MUX_BIT_9/s_top ), .ZN(n18197) );
  INV_X1 U17621 ( .A(\core_inst/MEM/MUX_LOAD/MUX_BIT_8/s_top ), .ZN(n18199) );
  INV_X1 U17622 ( .A(\core_inst/MEM/MUX_LOAD/MUX_BIT_10/s_top ), .ZN(n18225)
         );
  NOR3_X1 U17623 ( .A1(s_IFID_IR[26]), .A2(s_IFID_IR[30]), .A3(n14191), .ZN(
        n23282) );
  AOI221_X1 U17624 ( .B1(s_IFID_IR[22]), .B2(n19292), .C1(n19291), .C2(
        s_IFID_IR[25]), .A(n20045), .ZN(n20042) );
  OAI22_X1 U17625 ( .A1(s_IFID_IR[22]), .A2(n19292), .B1(s_IFID_IR[25]), .B2(
        n19291), .ZN(n20045) );
  NOR3_X1 U17626 ( .A1(net741458), .A2(net366531), .A3(n23283), .ZN(net712971)
         );
  NOR2_X1 U17627 ( .A1(net366211), .A2(net716215), .ZN(n23283) );
  NAND3_X1 U17628 ( .A1(n18179), .A2(n23284), .A3(n18135), .ZN(n18152) );
  AOI22_X1 U17629 ( .A1(n23285), .A2(net741565), .B1(n19282), .B2(n25745), 
        .ZN(n23284) );
  NAND2_X1 U17630 ( .A1(n26511), .A2(n18153), .ZN(n23285) );
  NAND2_X1 U17631 ( .A1(net741565), .A2(n26258), .ZN(net713425) );
  INV_X1 U17632 ( .A(n18152), .ZN(net713424) );
  AND2_X1 U17633 ( .A1(n20043), .A2(s_ID_rf_write_en), .ZN(n26270) );
  AOI221_X1 U17634 ( .B1(s_IFID_IR[24]), .B2(n19288), .C1(n19289), .C2(
        s_IFID_IR[23]), .A(n20044), .ZN(n20043) );
  OAI22_X1 U17635 ( .A1(s_IFID_IR[24]), .A2(n19288), .B1(s_IFID_IR[23]), .B2(
        n19289), .ZN(n20044) );
  OAI21_X1 U17636 ( .B1(n18175), .B2(n20133), .A(s_IFID_IR[30]), .ZN(n18158)
         );
  NOR3_X1 U17637 ( .A1(n14190), .A2(n18188), .A3(n20114), .ZN(n18181) );
  NAND3_X1 U17638 ( .A1(n14195), .A2(n18059), .A3(n24585), .ZN(n20114) );
  NOR3_X1 U17639 ( .A1(n14195), .A2(n18059), .A3(n20109), .ZN(n18146) );
  NAND2_X1 U17640 ( .A1(n20110), .A2(n14128), .ZN(n20109) );
  OAI21_X1 U17641 ( .B1(n18150), .B2(n20100), .A(n26777), .ZN(net713389) );
  OAI211_X1 U17642 ( .C1(n18062), .C2(n18170), .A(n18169), .B(n20105), .ZN(
        n20100) );
  INV_X1 U17643 ( .A(n18145), .ZN(n20105) );
  NAND2_X1 U17644 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[29] ), .ZN(
        n18205) );
  NAND2_X1 U17645 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[18] ), .ZN(
        n18216) );
  NAND2_X1 U17646 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[23] ), .ZN(
        n18211) );
  NAND2_X1 U17647 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[27] ), .ZN(
        n18207) );
  NAND2_X1 U17648 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[21] ), .ZN(
        n18213) );
  NAND2_X1 U17649 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[25] ), .ZN(
        n18209) );
  INV_X1 U17650 ( .A(\core_inst/MEM/MUX_LOAD/MUX_BIT_15/s_top ), .ZN(n18220)
         );
  NAND2_X1 U17651 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[16] ), .ZN(
        n18218) );
  NAND2_X1 U17652 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[31] ), .ZN(
        n18202) );
  NAND2_X1 U17653 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[26] ), .ZN(
        n18208) );
  NAND2_X1 U17654 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[30] ), .ZN(
        n18204) );
  NAND2_X1 U17655 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[20] ), .ZN(
        n18214) );
  NAND2_X1 U17656 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[24] ), .ZN(
        n18210) );
  NAND2_X1 U17657 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[17] ), .ZN(
        n18217) );
  NAND2_X1 U17658 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[22] ), .ZN(
        n18212) );
  NAND2_X1 U17659 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[19] ), .ZN(
        n18215) );
  NAND2_X1 U17660 ( .A1(n18203), .A2(\core_inst/s_DRAM_DLX_OUT[28] ), .ZN(
        n18206) );
  OAI211_X2 U17661 ( .C1(s_MEM_LOAD_TYPE[0]), .C2(n18219), .A(
        s_MEM_SIGNED_LOAD), .B(\core_inst/MEMWB_DATAOUT/DFF_15/N3 ), .ZN(
        n18201) );
  INV_X1 U17662 ( .A(n18198), .ZN(n18219) );
  NAND4_X1 U17663 ( .A1(s_IFID_IR[28]), .A2(s_IFID_IR[27]), .A3(s_IFID_IR[29]), 
        .A4(n20119), .ZN(n18179) );
  NOR3_X1 U17664 ( .A1(n14191), .A2(s_IFID_IR[26]), .A3(s_IFID_IR[30]), .ZN(
        n20119) );
  AND2_X1 U17665 ( .A1(n26274), .A2(n23286), .ZN(n26704) );
  NAND3_X1 U17666 ( .A1(n26270), .A2(n20041), .A3(n20042), .ZN(n23286) );
  NAND3_X1 U17667 ( .A1(net710387), .A2(net713389), .A3(n23287), .ZN(n26274)
         );
  OR2_X1 U17668 ( .A1(s_IFID_IR[30]), .A2(n26779), .ZN(n23287) );
  INV_X1 U17669 ( .A(net713439), .ZN(net713438) );
  OAI211_X1 U17670 ( .C1(n25769), .C2(n25768), .A(n23288), .B(n25767), .ZN(
        n25580) );
  NOR2_X1 U17671 ( .A1(n25765), .A2(n23026), .ZN(n23288) );
  INV_X1 U17672 ( .A(net712809), .ZN(net712808) );
  CLKBUF_X1 U17673 ( .A(net713454), .Z(net717696) );
  AOI21_X1 U17674 ( .B1(n24382), .B2(net717091), .A(n23289), .ZN(n24284) );
  CLKBUF_X1 U17675 ( .A(n24383), .Z(n23289) );
  CLKBUF_X1 U17676 ( .A(n25383), .Z(n23290) );
  CLKBUF_X1 U17677 ( .A(net713208), .Z(net742518) );
  NOR3_X1 U17678 ( .A1(net737706), .A2(n26533), .A3(n23291), .ZN(n26737) );
  AOI21_X1 U17679 ( .B1(n26532), .B2(n23292), .A(net729186), .ZN(n23291) );
  INV_X1 U17680 ( .A(n26531), .ZN(n23292) );
  AND3_X1 U17681 ( .A1(net780537), .A2(n23296), .A3(n23293), .ZN(n24787) );
  NAND2_X1 U17682 ( .A1(n23294), .A2(net732762), .ZN(n23293) );
  NAND3_X1 U17683 ( .A1(n23295), .A2(net712469), .A3(net750287), .ZN(n23294)
         );
  AND4_X1 U17684 ( .A1(net714487), .A2(net714486), .A3(net714488), .A4(
        net714489), .ZN(n23296) );
  CLKBUF_X1 U17685 ( .A(net738517), .Z(net738518) );
  CLKBUF_X1 U17686 ( .A(net733097), .Z(net755052) );
  CLKBUF_X1 U17687 ( .A(net713467), .Z(net749719) );
  INV_X1 U17688 ( .A(n23297), .ZN(n26571) );
  OAI21_X1 U17689 ( .B1(n26570), .B2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [24]), .A(net712838), .ZN(n23297) );
  INV_X1 U17690 ( .A(n23298), .ZN(n26736) );
  CLKBUF_X1 U17691 ( .A(net712473), .Z(net741975) );
  AOI21_X1 U17692 ( .B1(net713446), .B2(net717091), .A(n23299), .ZN(n26733) );
  BUF_X1 U17693 ( .A(n25512), .Z(n23299) );
  MUX2_X1 U17694 ( .A(net713892), .B(n26136), .S(net713606), .Z(net713910) );
  MUX2_X1 U17695 ( .A(net713728), .B(net713770), .S(net713606), .Z(net713993)
         );
  INV_X1 U17696 ( .A(n23300), .ZN(n25504) );
  OAI21_X1 U17697 ( .B1(n26214), .B2(n23301), .A(n26213), .ZN(n23300) );
  NAND2_X1 U17698 ( .A1(n24548), .A2(n23966), .ZN(n23301) );
  NOR2_X1 U17699 ( .A1(net712964), .A2(net760170), .ZN(n26740) );
  OAI21_X1 U17700 ( .B1(n23302), .B2(n26510), .A(net712971), .ZN(net712968) );
  XNOR2_X1 U17701 ( .A(n23303), .B(n26509), .ZN(n23302) );
  NAND2_X1 U17702 ( .A1(n26508), .A2(net712975), .ZN(n23303) );
  INV_X1 U17703 ( .A(net795273), .ZN(net712967) );
  NOR2_X1 U17704 ( .A1(net749894), .A2(n23304), .ZN(net714493) );
  NOR2_X1 U17705 ( .A1(n25999), .A2(net713726), .ZN(n23304) );
  NAND2_X1 U17706 ( .A1(n25999), .A2(net713736), .ZN(net714492) );
  OAI21_X1 U17707 ( .B1(net742087), .B2(net713892), .A(n26053), .ZN(net714228)
         );
  OAI22_X1 U17708 ( .A1(n26227), .A2(net767234), .B1(net713736), .B2(n26052), 
        .ZN(net714227) );
  CLKBUF_X1 U17709 ( .A(n26409), .Z(n23305) );
  AND2_X1 U17710 ( .A1(n24374), .A2(n23306), .ZN(n24199) );
  NOR2_X1 U17711 ( .A1(n24376), .A2(n24375), .ZN(n23306) );
  NAND2_X1 U17712 ( .A1(n25844), .A2(n23307), .ZN(n24565) );
  NOR2_X1 U17713 ( .A1(n23025), .A2(n25842), .ZN(n23307) );
  AOI21_X1 U17714 ( .B1(n25759), .B2(net717091), .A(n23308), .ZN(n25769) );
  NAND2_X1 U17715 ( .A1(n23309), .A2(net742483), .ZN(n23308) );
  MUX2_X1 U17716 ( .A(net713728), .B(net717087), .S(net717570), .Z(n23309) );
  NOR2_X1 U17717 ( .A1(net749894), .A2(n23310), .ZN(net713152) );
  OAI21_X1 U17718 ( .B1(net713554), .B2(net734121), .A(n23311), .ZN(n23310) );
  NAND2_X1 U17719 ( .A1(net713554), .A2(n26136), .ZN(n23311) );
  INV_X1 U17720 ( .A(net713892), .ZN(net734121) );
  OAI21_X1 U17721 ( .B1(n23312), .B2(n23313), .A(net713775), .ZN(n25767) );
  NOR2_X1 U17722 ( .A1(net762754), .A2(net762661), .ZN(n23313) );
  OAI22_X1 U17723 ( .A1(n24358), .A2(net717074), .B1(net728314), .B2(net748269), .ZN(n23312) );
  AOI22_X1 U17724 ( .A1(n24341), .A2(n23314), .B1(n24345), .B2(n23315), .ZN(
        n26221) );
  INV_X1 U17725 ( .A(n26200), .ZN(n23315) );
  INV_X1 U17726 ( .A(n23974), .ZN(n23314) );
  OAI21_X1 U17727 ( .B1(n23316), .B2(n23317), .A(net713863), .ZN(net713860) );
  OAI22_X1 U17728 ( .A1(net713773), .A2(net750287), .B1(net762753), .B2(
        net718355), .ZN(n23317) );
  OAI222_X1 U17729 ( .A1(net717055), .A2(net713810), .B1(n24357), .B2(
        net767206), .C1(net717074), .C2(net755699), .ZN(n23316) );
  AOI22_X1 U17730 ( .A1(net713869), .A2(net713779), .B1(net713870), .B2(
        net767211), .ZN(net713859) );
  AOI22_X1 U17731 ( .A1(net713785), .A2(n26137), .B1(net713873), .B2(net713874), .ZN(net713858) );
  OAI22_X1 U17732 ( .A1(net767206), .A2(net717074), .B1(n24357), .B2(net713810), .ZN(net714491) );
  OAI22_X1 U17733 ( .A1(net713773), .A2(net717055), .B1(net762754), .B2(
        net755699), .ZN(net714490) );
  NAND2_X1 U17734 ( .A1(net714965), .A2(net715241), .ZN(n25859) );
  AOI21_X1 U17735 ( .B1(n26177), .B2(n23318), .A(n23319), .ZN(n25408) );
  NAND2_X1 U17736 ( .A1(n23320), .A2(net718367), .ZN(n23319) );
  MUX2_X1 U17737 ( .A(net713770), .B(n23322), .S(net749732), .Z(n23320) );
  AND2_X1 U17738 ( .A1(net713154), .A2(n25662), .ZN(n23322) );
  NOR2_X1 U17739 ( .A1(n26175), .A2(n23321), .ZN(n23318) );
  AND2_X1 U17740 ( .A1(n24177), .A2(n25413), .ZN(n23321) );
  NOR2_X1 U17741 ( .A1(n23324), .A2(n23323), .ZN(n25428) );
  NOR2_X1 U17742 ( .A1(n24192), .A2(net742304), .ZN(n23324) );
  AND2_X1 U17743 ( .A1(n23325), .A2(n25831), .ZN(n24285) );
  NOR2_X1 U17744 ( .A1(n25830), .A2(n25829), .ZN(n23325) );
  NOR2_X1 U17745 ( .A1(n24027), .A2(n25849), .ZN(n23326) );
  AND3_X1 U17746 ( .A1(n23326), .A2(n26048), .A3(n26049), .ZN(n26223) );
  NAND3_X1 U17747 ( .A1(n23327), .A2(n23328), .A3(net717091), .ZN(n26606) );
  OAI21_X1 U17748 ( .B1(n23333), .B2(net714858), .A(n23329), .ZN(n23328) );
  NOR2_X1 U17749 ( .A1(n24538), .A2(net780578), .ZN(n23329) );
  OR3_X1 U17750 ( .A1(n24286), .A2(n24818), .A3(n24292), .ZN(n23333) );
  OAI211_X1 U17751 ( .C1(net715200), .C2(n23332), .A(n23330), .B(n24352), .ZN(
        n23327) );
  XNOR2_X1 U17752 ( .A(n23331), .B(n26064), .ZN(n23330) );
  XOR2_X1 U17753 ( .A(n24531), .B(net716221), .Z(n23331) );
  NOR3_X1 U17754 ( .A1(n24286), .A2(n24818), .A3(n24292), .ZN(n23332) );
  OAI22_X1 U17755 ( .A1(net767205), .A2(n4344), .B1(net718134), .B2(n24815), 
        .ZN(n23334) );
  NOR2_X1 U17756 ( .A1(net762680), .A2(n4343), .ZN(n23335) );
  NOR2_X1 U17757 ( .A1(n23334), .A2(n23335), .ZN(n23336) );
  NAND2_X1 U17758 ( .A1(net742331), .A2(n17957), .ZN(n23337) );
  NAND3_X1 U17759 ( .A1(n23336), .A2(n23337), .A3(n25760), .ZN(n26143) );
  AND3_X1 U17760 ( .A1(n24290), .A2(net749930), .A3(n23338), .ZN(n24818) );
  OR2_X1 U17761 ( .A1(n23968), .A2(n23339), .ZN(n23338) );
  CLKBUF_X1 U17762 ( .A(n25825), .Z(n23339) );
  NAND3_X1 U17763 ( .A1(n23340), .A2(n25386), .A3(n25385), .ZN(n24531) );
  AOI21_X1 U17764 ( .B1(n24193), .B2(net365821), .A(n23341), .ZN(n23340) );
  CLKBUF_X1 U17765 ( .A(n25387), .Z(n23341) );
  AND2_X1 U17766 ( .A1(n23342), .A2(n26192), .ZN(n26251) );
  NAND3_X1 U17767 ( .A1(n26191), .A2(n24301), .A3(n26194), .ZN(n23342) );
  OAI22_X1 U17768 ( .A1(n23343), .A2(n23344), .B1(net742087), .B2(net713767), 
        .ZN(n26567) );
  NOR2_X1 U17769 ( .A1(n23345), .A2(net742436), .ZN(n23344) );
  INV_X1 U17770 ( .A(net796212), .ZN(net742436) );
  OAI21_X1 U17771 ( .B1(n23345), .B2(net734022), .A(net713863), .ZN(n23343) );
  NOR2_X1 U17772 ( .A1(net762753), .A2(net713810), .ZN(n23345) );
  NOR2_X1 U17773 ( .A1(n26058), .A2(net742243), .ZN(n23346) );
  AOI21_X1 U17774 ( .B1(n23347), .B2(net717091), .A(n23348), .ZN(n25768) );
  NAND3_X1 U17775 ( .A1(n25381), .A2(net714194), .A3(n23349), .ZN(n23348) );
  MUX2_X1 U17776 ( .A(net713726), .B(n25662), .S(net717570), .Z(n23349) );
  INV_X1 U17777 ( .A(n25759), .ZN(n23347) );
  XNOR2_X1 U17778 ( .A(n23350), .B(n23351), .ZN(n25759) );
  INV_X1 U17779 ( .A(n23353), .ZN(n23351) );
  CLKBUF_X1 U17780 ( .A(n24281), .Z(n23353) );
  NOR2_X1 U17781 ( .A1(n23968), .A2(n23352), .ZN(n23350) );
  NOR2_X1 U17782 ( .A1(n24551), .A2(n25513), .ZN(n23352) );
  AND2_X1 U17783 ( .A1(n26227), .A2(n23354), .ZN(n26225) );
  AND2_X1 U17784 ( .A1(net713564), .A2(n26228), .ZN(n23354) );
  NAND2_X1 U17785 ( .A1(net717789), .A2(n522), .ZN(n23355) );
  OAI221_X1 U17786 ( .B1(net749972), .B2(n1716), .C1(net750086), .C2(n4358), 
        .A(n23355), .ZN(n23356) );
  AOI221_X1 U17787 ( .B1(n24295), .B2(n17674), .C1(net749806), .C2(n25332), 
        .A(n23356), .ZN(n23357) );
  INV_X1 U17788 ( .A(n23357), .ZN(n26001) );
  XNOR2_X1 U17789 ( .A(n23358), .B(
        \core_inst/IF_stage/PLUS4_ADDER/RES_GENERATOR/CSA_15/sum_rca_0[1] ), 
        .ZN(n25446) );
  OR2_X1 U17790 ( .A1(n23359), .A2(net712847), .ZN(n23358) );
  NAND2_X1 U17791 ( .A1(
        \core_inst/IF_stage/PLUS4_ADDER/RES_GENERATOR/CSA_15/RCA_1/cout_tmp[0] ), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [29]), .ZN(n23359) );
  NOR2_X1 U17792 ( .A1(n24548), .A2(net749534), .ZN(n23360) );
  NOR2_X1 U17793 ( .A1(n23361), .A2(net713154), .ZN(net713442) );
  XNOR2_X1 U17794 ( .A(n23362), .B(n23363), .ZN(n23361) );
  NOR2_X1 U17795 ( .A1(n25971), .A2(n24344), .ZN(n23363) );
  NAND2_X1 U17796 ( .A1(n23364), .A2(n26020), .ZN(n23362) );
  NAND3_X1 U17797 ( .A1(n25424), .A2(n23365), .A3(net740526), .ZN(n23364) );
  NOR2_X1 U17798 ( .A1(net714631), .A2(n24568), .ZN(n23365) );
  INV_X1 U17799 ( .A(net739130), .ZN(net714631) );
  OAI22_X1 U17800 ( .A1(n23366), .A2(n23367), .B1(n26046), .B2(n25946), .ZN(
        n25947) );
  NAND2_X1 U17801 ( .A1(n26025), .A2(n26024), .ZN(n23367) );
  NAND3_X1 U17802 ( .A1(n26026), .A2(n22812), .A3(n24536), .ZN(n23366) );
  INV_X1 U17803 ( .A(net767221), .ZN(net778669) );
  NOR2_X1 U17804 ( .A1(n25579), .A2(net778669), .ZN(n23368) );
  NAND2_X1 U17805 ( .A1(net733229), .A2(net749427), .ZN(net733227) );
  OAI211_X1 U17806 ( .C1(n26223), .C2(n24278), .A(n23369), .B(n26221), .ZN(
        n26247) );
  AND4_X1 U17807 ( .A1(n26202), .A2(n26211), .A3(n26207), .A4(n26206), .ZN(
        n23369) );
  NAND2_X1 U17808 ( .A1(net724352), .A2(net741531), .ZN(net724354) );
  NAND2_X1 U17809 ( .A1(net716215), .A2(n23370), .ZN(net724353) );
  NAND2_X1 U17810 ( .A1(net741282), .A2(net741531), .ZN(n23370) );
  AOI21_X1 U17811 ( .B1(n23371), .B2(n22830), .A(n23372), .ZN(net724352) );
  NAND2_X1 U17812 ( .A1(n24563), .A2(n23373), .ZN(n23372) );
  INV_X1 U17813 ( .A(n26238), .ZN(n23373) );
  NAND3_X1 U17814 ( .A1(n26252), .A2(n26251), .A3(n25504), .ZN(n23371) );
  NAND2_X1 U17815 ( .A1(n26232), .A2(n23374), .ZN(n26244) );
  OAI21_X1 U17816 ( .B1(n26228), .B2(net713564), .A(n26227), .ZN(n23374) );
  NOR2_X1 U17817 ( .A1(n4346), .A2(net741959), .ZN(n23375) );
  AOI21_X1 U17818 ( .B1(n24295), .B2(n25345), .A(n23375), .ZN(n23376) );
  NOR2_X1 U17819 ( .A1(net749972), .A2(n1752), .ZN(n23377) );
  AOI221_X1 U17820 ( .B1(net717789), .B2(net741582), .C1(net749806), .C2(
        n17670), .A(n23377), .ZN(n23378) );
  NAND2_X1 U17821 ( .A1(n23376), .A2(n23378), .ZN(n26168) );
  NAND2_X1 U17822 ( .A1(n23379), .A2(n26230), .ZN(n26243) );
  NAND3_X1 U17823 ( .A1(n26229), .A2(net742507), .A3(net713561), .ZN(n23379)
         );
  NAND4_X1 U17824 ( .A1(n26245), .A2(n26244), .A3(n23380), .A4(n26242), .ZN(
        n26238) );
  NAND3_X1 U17825 ( .A1(n26232), .A2(n23381), .A3(n26243), .ZN(n23380) );
  NAND3_X1 U17826 ( .A1(n23382), .A2(n23383), .A3(n23384), .ZN(n25396) );
  AOI22_X1 U17827 ( .A1(n26211), .A2(n23385), .B1(net755740), .B2(n26210), 
        .ZN(n23384) );
  NOR2_X1 U17828 ( .A1(n24196), .A2(n26208), .ZN(n23385) );
  AOI21_X1 U17829 ( .B1(net713606), .B2(net713607), .A(n23386), .ZN(n23383) );
  INV_X1 U17830 ( .A(n26229), .ZN(n23386) );
  NAND4_X1 U17831 ( .A1(n23387), .A2(n26211), .A3(n26207), .A4(n26206), .ZN(
        n23382) );
  OAI22_X1 U17832 ( .A1(net750238), .A2(n24293), .B1(net713614), .B2(n24198), 
        .ZN(n23387) );
  NAND3_X1 U17833 ( .A1(n23390), .A2(n23389), .A3(n23388), .ZN(n26107) );
  OR2_X1 U17834 ( .A1(net742413), .A2(n1730), .ZN(n23388) );
  OR2_X1 U17835 ( .A1(net742223), .A2(n4356), .ZN(n23389) );
  AOI22_X1 U17836 ( .A1(net718341), .A2(n24604), .B1(n24275), .B2(n25351), 
        .ZN(n23390) );
  NAND2_X1 U17837 ( .A1(n23391), .A2(n23392), .ZN(n26052) );
  NOR2_X1 U17838 ( .A1(n23393), .A2(n23394), .ZN(n23392) );
  NOR2_X1 U17839 ( .A1(net741959), .A2(n4355), .ZN(n23394) );
  OAI22_X1 U17840 ( .A1(net749972), .A2(n1730), .B1(net749495), .B2(n4356), 
        .ZN(n23393) );
  AOI22_X1 U17841 ( .A1(net742331), .A2(n25333), .B1(n24295), .B2(n17675), 
        .ZN(n23391) );
  NAND2_X1 U17842 ( .A1(n23395), .A2(net717091), .ZN(n26580) );
  XNOR2_X1 U17843 ( .A(n23397), .B(n23396), .ZN(n23395) );
  XNOR2_X1 U17844 ( .A(n24571), .B(net714729), .ZN(n23396) );
  INV_X1 U17845 ( .A(net713612), .ZN(net714729) );
  AOI21_X1 U17846 ( .B1(n25939), .B2(net742423), .A(n25373), .ZN(n23397) );
  NAND3_X1 U17847 ( .A1(n24332), .A2(net758644), .A3(n25503), .ZN(n23398) );
  NAND2_X1 U17848 ( .A1(n24292), .A2(net758644), .ZN(n23399) );
  NAND3_X1 U17849 ( .A1(n23398), .A2(n23399), .A3(net778368), .ZN(net713168)
         );
  NOR2_X1 U17850 ( .A1(n23400), .A2(n23401), .ZN(n26163) );
  OAI21_X1 U17851 ( .B1(net713564), .B2(net714871), .A(net714877), .ZN(n23401)
         );
  OAI211_X1 U17852 ( .C1(n25986), .C2(net742092), .A(n23402), .B(n23403), .ZN(
        n23400) );
  NAND2_X1 U17853 ( .A1(n24322), .A2(net750274), .ZN(n23403) );
  NAND2_X1 U17854 ( .A1(net750025), .A2(net713753), .ZN(n23402) );
  INV_X1 U17855 ( .A(net755040), .ZN(net750290) );
  AOI21_X1 U17856 ( .B1(n23404), .B2(n23948), .A(n25394), .ZN(net755040) );
  NOR2_X1 U17857 ( .A1(n24265), .A2(n24029), .ZN(n23404) );
  NOR2_X1 U17858 ( .A1(n23405), .A2(n23406), .ZN(n25466) );
  NOR2_X1 U17859 ( .A1(net750090), .A2(net742304), .ZN(n23406) );
  NOR2_X1 U17860 ( .A1(n24548), .A2(net796014), .ZN(n23405) );
  NAND4_X1 U17861 ( .A1(n23407), .A2(n23408), .A3(n23409), .A4(n23410), .ZN(
        n26175) );
  NAND2_X1 U17862 ( .A1(net713748), .A2(net749387), .ZN(n23410) );
  AOI21_X1 U17863 ( .B1(net737713), .B2(net748269), .A(net713751), .ZN(n23409)
         );
  NAND2_X1 U17864 ( .A1(n24355), .A2(net749812), .ZN(n23408) );
  NAND2_X1 U17865 ( .A1(net712468), .A2(net713754), .ZN(n23407) );
  XNOR2_X1 U17866 ( .A(n23411), .B(net716215), .ZN(n24178) );
  NAND2_X1 U17867 ( .A1(n23976), .A2(n25822), .ZN(n23411) );
  NOR2_X1 U17868 ( .A1(net713854), .A2(n23412), .ZN(net712462) );
  OR2_X1 U17869 ( .A1(n24203), .A2(n24550), .ZN(n23412) );
  INV_X1 U17870 ( .A(net713857), .ZN(net713854) );
  OR2_X1 U17871 ( .A1(net717510), .A2(n23413), .ZN(n25789) );
  NAND2_X1 U17872 ( .A1(n24206), .A2(n26143), .ZN(n23413) );
  OAI21_X1 U17873 ( .B1(n25407), .B2(n25408), .A(n23414), .ZN(net760170) );
  AND2_X1 U17874 ( .A1(n25409), .A2(n25410), .ZN(n23414) );
  OAI211_X1 U17875 ( .C1(n25407), .C2(n25408), .A(n25409), .B(n25410), .ZN(
        net712965) );
  NAND4_X1 U17876 ( .A1(n23415), .A2(n23416), .A3(n23417), .A4(n23418), .ZN(
        n26174) );
  NAND2_X1 U17877 ( .A1(net749500), .A2(net717875), .ZN(n23418) );
  NAND2_X1 U17878 ( .A1(net749898), .A2(net749260), .ZN(n23417) );
  AOI22_X1 U17879 ( .A1(n24577), .A2(net750158), .B1(n24272), .B2(net755238), 
        .ZN(n23416) );
  NAND2_X1 U17880 ( .A1(n24330), .A2(net749534), .ZN(n23415) );
  AOI21_X1 U17881 ( .B1(n23422), .B2(n26176), .A(n23419), .ZN(n25407) );
  NAND2_X1 U17882 ( .A1(n23420), .A2(net739078), .ZN(n23419) );
  MUX2_X1 U17883 ( .A(n23423), .B(net713726), .S(net749732), .Z(n23420) );
  AND2_X1 U17884 ( .A1(net713154), .A2(net713728), .ZN(n23423) );
  AND2_X1 U17885 ( .A1(n23421), .A2(n26178), .ZN(n23422) );
  INV_X1 U17886 ( .A(n26174), .ZN(n23421) );
  NAND2_X1 U17887 ( .A1(n26189), .A2(n23424), .ZN(n26220) );
  AOI21_X1 U17888 ( .B1(net749823), .B2(n23426), .A(n23425), .ZN(n23424) );
  NOR2_X1 U17889 ( .A1(n24274), .A2(n24318), .ZN(n23425) );
  INV_X1 U17890 ( .A(n26188), .ZN(n23426) );
  AOI21_X1 U17891 ( .B1(n23428), .B2(n23429), .A(n23427), .ZN(n25395) );
  NAND4_X1 U17892 ( .A1(n26202), .A2(n26211), .A3(n26207), .A4(n26206), .ZN(
        n23427) );
  NAND2_X1 U17893 ( .A1(n24543), .A2(n26200), .ZN(n23429) );
  AOI22_X1 U17894 ( .A1(n23430), .A2(n26221), .B1(n26199), .B2(net713633), 
        .ZN(n23428) );
  OAI21_X1 U17895 ( .B1(n24544), .B2(n23431), .A(n26196), .ZN(n23430) );
  INV_X1 U17896 ( .A(n26223), .ZN(n23431) );
  NOR3_X1 U17897 ( .A1(n25395), .A2(n26241), .A3(n25396), .ZN(n24563) );
  NOR3_X2 U17898 ( .A1(n26203), .A2(n23432), .A3(n26233), .ZN(n26232) );
  AND2_X1 U17899 ( .A1(net713151), .A2(net713554), .ZN(n23432) );
  OAI211_X1 U17900 ( .C1(n26226), .C2(n23433), .A(n26232), .B(n23434), .ZN(
        n26245) );
  INV_X1 U17901 ( .A(n26225), .ZN(n23434) );
  NOR3_X1 U17902 ( .A1(net746701), .A2(n26224), .A3(net762674), .ZN(n23433) );
  NOR2_X1 U17903 ( .A1(n26408), .A2(net713151), .ZN(net715351) );
  NAND2_X1 U17904 ( .A1(net712467), .A2(n23435), .ZN(net713148) );
  AND2_X1 U17905 ( .A1(net734022), .A2(net713863), .ZN(n23435) );
  NAND2_X1 U17906 ( .A1(n23436), .A2(net713570), .ZN(net714544) );
  XNOR2_X1 U17907 ( .A(net713934), .B(net716215), .ZN(n23436) );
  INV_X1 U17908 ( .A(n23437), .ZN(n25848) );
  OAI22_X1 U17909 ( .A1(net718133), .A2(n23268), .B1(net749926), .B2(n680), 
        .ZN(n23437) );
  OR2_X1 U17910 ( .A1(n23438), .A2(n23439), .ZN(n25338) );
  MUX2_X1 U17911 ( .A(n23440), .B(n23441), .S(net742315), .Z(n23439) );
  MUX2_X1 U17912 ( .A(net767234), .B(net713736), .S(n26200), .Z(n23441) );
  NAND2_X1 U17913 ( .A1(net713767), .A2(n23442), .ZN(n23440) );
  MUX2_X1 U17914 ( .A(net713726), .B(n25662), .S(n26200), .Z(n23442) );
  MUX2_X1 U17915 ( .A(n25947), .B(net714378), .S(net718367), .Z(n23438) );
  XNOR2_X1 U17916 ( .A(n23443), .B(n23444), .ZN(n24235) );
  AND2_X1 U17917 ( .A1(n24352), .A2(net755105), .ZN(n23444) );
  INV_X1 U17918 ( .A(net715200), .ZN(net755105) );
  NOR3_X1 U17919 ( .A1(n24286), .A2(n24818), .A3(n24292), .ZN(n23443) );
  AOI22_X1 U17920 ( .A1(n24306), .A2(net767211), .B1(net713870), .B2(net713779), .ZN(net778055) );
  NAND2_X1 U17921 ( .A1(n26163), .A2(net713785), .ZN(net778056) );
  AOI22_X1 U17922 ( .A1(n26050), .A2(net713874), .B1(n26203), .B2(n26136), 
        .ZN(net778057) );
  NOR2_X1 U17923 ( .A1(net762680), .A2(n4367), .ZN(n23445) );
  OAI22_X1 U17924 ( .A1(net717106), .A2(n1738), .B1(net718361), .B2(n4368), 
        .ZN(n23446) );
  NOR2_X1 U17925 ( .A1(n23445), .A2(n23446), .ZN(n23447) );
  AOI22_X1 U17926 ( .A1(n24295), .A2(n14464), .B1(net780566), .B2(n25331), 
        .ZN(n23448) );
  NAND2_X1 U17927 ( .A1(n23447), .A2(n23448), .ZN(n25991) );
  AOI21_X1 U17928 ( .B1(n24295), .B2(n17663), .A(n23449), .ZN(n25827) );
  NOR2_X1 U17929 ( .A1(n23450), .A2(n23451), .ZN(n26101) );
  OAI22_X1 U17930 ( .A1(n1724), .A2(net715419), .B1(n25311), .B2(net742223), 
        .ZN(n23451) );
  OAI22_X1 U17931 ( .A1(n25391), .A2(n25363), .B1(net715422), .B2(n4373), .ZN(
        n23450) );
  NOR2_X1 U17932 ( .A1(n23452), .A2(n23453), .ZN(n25851) );
  OAI22_X1 U17933 ( .A1(net765744), .A2(n1718), .B1(net749495), .B2(n25308), 
        .ZN(n23453) );
  NOR2_X1 U17934 ( .A1(net718133), .A2(n23267), .ZN(n23452) );
  OAI22_X1 U17935 ( .A1(net767340), .A2(n23269), .B1(net717615), .B2(n22676), 
        .ZN(n23454) );
  NAND2_X1 U17936 ( .A1(n24320), .A2(n25330), .ZN(n23455) );
  OAI221_X1 U17937 ( .B1(net749495), .B2(n25283), .C1(net765744), .C2(n1722), 
        .A(n23455), .ZN(n23456) );
  OR2_X1 U17938 ( .A1(n23454), .A2(n23456), .ZN(n26197) );
  AOI21_X1 U17939 ( .B1(n23457), .B2(net713813), .A(n22829), .ZN(net714106) );
  NOR2_X1 U17940 ( .A1(n25598), .A2(net749454), .ZN(n23457) );
  INV_X1 U17941 ( .A(n23458), .ZN(n26064) );
  MUX2_X1 U17942 ( .A(n17924), .B(n25392), .S(net787518), .Z(n23458) );
  NAND2_X1 U17943 ( .A1(n23459), .A2(n23460), .ZN(n26046) );
  AOI22_X1 U17944 ( .A1(net742157), .A2(n26148), .B1(net767207), .B2(net714249), .ZN(n23459) );
  INV_X1 U17945 ( .A(n23461), .ZN(n25850) );
  OAI22_X1 U17946 ( .A1(n4388), .A2(net762680), .B1(n874), .B2(net765629), 
        .ZN(n23461) );
  NAND3_X1 U17947 ( .A1(n23462), .A2(n23463), .A3(n23464), .ZN(n26085) );
  NAND2_X1 U17948 ( .A1(n24275), .A2(n25343), .ZN(n23464) );
  NAND2_X1 U17949 ( .A1(net750031), .A2(n25328), .ZN(n23463) );
  AOI22_X1 U17950 ( .A1(net742412), .A2(\core_inst/MEMWB_ALUOUT/DFF_30/N3 ), 
        .B1(net750111), .B2(n482), .ZN(n23462) );
  NAND2_X1 U17951 ( .A1(net796255), .A2(n23465), .ZN(n26672) );
  INV_X1 U17952 ( .A(n23466), .ZN(n23465) );
  OAI21_X1 U17953 ( .B1(n26575), .B2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [10]), .A(n26459), .ZN(n23466) );
  OAI21_X1 U17954 ( .B1(n26579), .B2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [16]), .A(n26578), .ZN(n23467) );
  OR3_X1 U17955 ( .A1(n23469), .A2(n23470), .A3(n23471), .ZN(n25885) );
  NOR2_X1 U17956 ( .A1(net749679), .A2(net746701), .ZN(n23471) );
  NOR2_X1 U17957 ( .A1(net755683), .A2(n24543), .ZN(n23470) );
  NOR2_X1 U17958 ( .A1(net713151), .A2(n23468), .ZN(n23469) );
  INV_X1 U17959 ( .A(n24321), .ZN(n23468) );
  MUX2_X1 U17960 ( .A(n23472), .B(n23473), .S(net749306), .Z(net714356) );
  MUX2_X1 U17961 ( .A(net713728), .B(net713770), .S(n24171), .Z(n23473) );
  NAND2_X1 U17962 ( .A1(n24091), .A2(net713892), .ZN(n23472) );
  NAND2_X1 U17963 ( .A1(n26028), .A2(net714275), .ZN(net714355) );
  NOR2_X1 U17964 ( .A1(n23474), .A2(n23475), .ZN(n25847) );
  AND2_X1 U17965 ( .A1(n24320), .A2(n25317), .ZN(n23475) );
  OAI22_X1 U17966 ( .A1(net749972), .A2(n1740), .B1(net749495), .B2(n25312), 
        .ZN(n23474) );
  NOR2_X1 U17967 ( .A1(net715172), .A2(net715171), .ZN(net715170) );
  OAI222_X1 U17968 ( .A1(net741959), .A2(n25282), .B1(net765744), .B2(n1736), 
        .C1(net749495), .C2(net740721), .ZN(n23476) );
  OAI22_X1 U17969 ( .A1(net718133), .A2(n23270), .B1(net715058), .B2(n25320), 
        .ZN(n23477) );
  OR2_X2 U17970 ( .A1(n23476), .A2(n23477), .ZN(n26208) );
  NAND2_X1 U17971 ( .A1(n23478), .A2(n23479), .ZN(net714378) );
  NAND4_X1 U17972 ( .A1(n25421), .A2(n25466), .A3(n22812), .A4(n26027), .ZN(
        n23479) );
  NAND4_X1 U17973 ( .A1(n25959), .A2(n25989), .A3(n25428), .A4(n24536), .ZN(
        n23478) );
  NAND2_X1 U17974 ( .A1(n24193), .A2(n25328), .ZN(n23480) );
  OAI21_X1 U17975 ( .B1(net749972), .B2(n1734), .A(n23480), .ZN(n23481) );
  OAI222_X1 U17976 ( .A1(net718133), .A2(n22688), .B1(net765629), .B2(n22672), 
        .C1(net780584), .C2(n25349), .ZN(n23482) );
  NOR2_X2 U17977 ( .A1(n23481), .A2(n23482), .ZN(net713554) );
  NOR2_X1 U17978 ( .A1(n23483), .A2(n23484), .ZN(n25826) );
  NOR2_X1 U17979 ( .A1(n4337), .A2(n25595), .ZN(n23484) );
  OAI22_X1 U17980 ( .A1(net717106), .A2(n1706), .B1(net718361), .B2(n25346), 
        .ZN(n23483) );
  NAND3_X1 U17981 ( .A1(n26158), .A2(net714873), .A3(n23485), .ZN(n25886) );
  NAND2_X1 U17982 ( .A1(net749489), .A2(n25909), .ZN(n23485) );
  NOR2_X1 U17983 ( .A1(n26225), .A2(n23486), .ZN(n26231) );
  NAND2_X1 U17984 ( .A1(n23487), .A2(n23488), .ZN(n23486) );
  INV_X1 U17985 ( .A(n26224), .ZN(n23488) );
  NAND3_X1 U17986 ( .A1(net742473), .A2(net762674), .A3(n24326), .ZN(n23487)
         );
  INV_X1 U17987 ( .A(n23489), .ZN(n25854) );
  OAI22_X1 U17988 ( .A1(n23263), .A2(net767341), .B1(net742037), .B2(n22675), 
        .ZN(n23489) );
  NOR2_X1 U17989 ( .A1(n23490), .A2(n23491), .ZN(n25839) );
  OAI22_X1 U17990 ( .A1(net749972), .A2(n1710), .B1(net714943), .B2(n4401), 
        .ZN(n23491) );
  NOR2_X1 U17991 ( .A1(n25358), .A2(net767340), .ZN(n23490) );
  OAI211_X1 U17992 ( .C1(n26163), .C2(net739078), .A(n25989), .B(n23492), .ZN(
        n26407) );
  NAND2_X1 U17993 ( .A1(n25996), .A2(net739078), .ZN(n23492) );
  NAND2_X1 U17994 ( .A1(net742612), .A2(n23493), .ZN(n26711) );
  INV_X1 U17995 ( .A(n23494), .ZN(n23493) );
  OAI21_X1 U17996 ( .B1(n26457), .B2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [26]), .A(n26558), .ZN(n23494) );
  INV_X1 U17997 ( .A(net713614), .ZN(net714394) );
  MUX2_X1 U17998 ( .A(n26088), .B(n5587), .S(net741686), .Z(net713614) );
  OAI22_X1 U17999 ( .A1(net718336), .A2(n25308), .B1(net718432), .B2(n1718), 
        .ZN(net765677) );
  MUX2_X1 U18000 ( .A(n25986), .B(n23495), .S(net750176), .Z(net713873) );
  INV_X1 U18001 ( .A(n25985), .ZN(n23495) );
  NOR2_X1 U18002 ( .A1(n23496), .A2(n23497), .ZN(n25986) );
  OAI22_X1 U18003 ( .A1(n24278), .A2(n25781), .B1(net755134), .B2(n25782), 
        .ZN(n23497) );
  OAI22_X1 U18004 ( .A1(n24558), .A2(net749732), .B1(net713607), .B2(n22836), 
        .ZN(n23496) );
  AOI22_X1 U18005 ( .A1(net750238), .A2(net749967), .B1(net750158), .B2(n24311), .ZN(n25762) );
  INV_X1 U18006 ( .A(net715173), .ZN(net715169) );
  OAI22_X1 U18007 ( .A1(n1677), .A2(net767341), .B1(net715058), .B2(n25322), 
        .ZN(net715173) );
  NAND2_X1 U18008 ( .A1(n26249), .A2(n23498), .ZN(n26254) );
  NAND2_X1 U18009 ( .A1(n26246), .A2(n23499), .ZN(n23498) );
  INV_X1 U18010 ( .A(n26247), .ZN(n23499) );
  NAND3_X1 U18011 ( .A1(n23500), .A2(n22830), .A3(n26254), .ZN(n26508) );
  OAI21_X1 U18012 ( .B1(n26252), .B2(n23501), .A(n26251), .ZN(n23500) );
  INV_X1 U18013 ( .A(n26250), .ZN(n23501) );
  NAND2_X1 U18014 ( .A1(n23502), .A2(n23503), .ZN(n26246) );
  NAND3_X1 U18015 ( .A1(n23504), .A2(n26245), .A3(n26244), .ZN(n23503) );
  NOR2_X1 U18016 ( .A1(n22847), .A2(n26243), .ZN(n23504) );
  NAND4_X1 U18017 ( .A1(n26241), .A2(n26244), .A3(n23505), .A4(n26240), .ZN(
        n23502) );
  INV_X1 U18018 ( .A(n26239), .ZN(n23505) );
  AND2_X2 U18019 ( .A1(n26561), .A2(n23506), .ZN(n25366) );
  NAND2_X1 U18020 ( .A1(n25515), .A2(n24094), .ZN(n23506) );
  NAND4_X1 U18021 ( .A1(n23507), .A2(n23508), .A3(n23509), .A4(n23510), .ZN(
        n25750) );
  XOR2_X1 U18022 ( .A(net342954), .B(n1637), .Z(n23510) );
  XOR2_X1 U18023 ( .A(n25590), .B(n5181), .Z(n23509) );
  XNOR2_X1 U18024 ( .A(n25592), .B(n1643), .ZN(n23508) );
  NOR2_X1 U18025 ( .A1(n23511), .A2(n23512), .ZN(n23507) );
  XNOR2_X1 U18026 ( .A(net342961), .B(n5607), .ZN(n23512) );
  XNOR2_X1 U18027 ( .A(net366410), .B(n1641), .ZN(n23511) );
  NAND2_X1 U18028 ( .A1(net755708), .A2(n23513), .ZN(net712737) );
  AOI21_X1 U18029 ( .B1(n5576), .B2(n26671), .A(n26572), .ZN(n23513) );
  NAND3_X1 U18030 ( .A1(n23516), .A2(n23515), .A3(n23514), .ZN(n26087) );
  OR2_X1 U18031 ( .A1(net718337), .A2(n4368), .ZN(n23514) );
  OR2_X1 U18032 ( .A1(net742413), .A2(n1738), .ZN(n23515) );
  AOI22_X1 U18033 ( .A1(net718341), .A2(n24603), .B1(n24275), .B2(n25353), 
        .ZN(n23516) );
  NAND2_X2 U18034 ( .A1(n23517), .A2(n23518), .ZN(net714559) );
  OR2_X1 U18035 ( .A1(net716237), .A2(net81266), .ZN(n23518) );
  NAND2_X1 U18036 ( .A1(n26087), .A2(net716237), .ZN(n23517) );
  NAND3_X1 U18037 ( .A1(net712975), .A2(n26508), .A3(n23519), .ZN(net713496)
         );
  NOR2_X1 U18038 ( .A1(n23520), .A2(n26510), .ZN(n23519) );
  NAND2_X1 U18039 ( .A1(n23520), .A2(n26255), .ZN(net713495) );
  INV_X1 U18040 ( .A(n26509), .ZN(n23520) );
  NAND2_X1 U18041 ( .A1(n26254), .A2(n23521), .ZN(net712975) );
  NAND3_X1 U18042 ( .A1(n26248), .A2(n25504), .A3(n26249), .ZN(n23521) );
  INV_X1 U18043 ( .A(n23522), .ZN(n26132) );
  AOI21_X1 U18044 ( .B1(n25898), .B2(n23977), .A(net714861), .ZN(n23522) );
  NAND2_X1 U18045 ( .A1(n23528), .A2(n23529), .ZN(net729530) );
  NAND2_X1 U18046 ( .A1(n25424), .A2(n23531), .ZN(n23529) );
  AND2_X1 U18047 ( .A1(n26020), .A2(n23532), .ZN(n23528) );
  AND2_X1 U18048 ( .A1(n23533), .A2(n23534), .ZN(n23532) );
  AOI21_X1 U18049 ( .B1(n23524), .B2(n23523), .A(n23527), .ZN(net725022) );
  OAI21_X1 U18050 ( .B1(n23525), .B2(n26021), .A(net717091), .ZN(n23527) );
  NAND2_X1 U18051 ( .A1(n26020), .A2(n23533), .ZN(n23524) );
  INV_X1 U18052 ( .A(n25971), .ZN(n23533) );
  NAND2_X1 U18053 ( .A1(n23530), .A2(n23523), .ZN(net729531) );
  NOR2_X1 U18054 ( .A1(n23534), .A2(n24344), .ZN(n23523) );
  INV_X1 U18055 ( .A(n23525), .ZN(n23534) );
  XNOR2_X1 U18056 ( .A(n24296), .B(net713633), .ZN(n23525) );
  AND2_X1 U18057 ( .A1(n25424), .A2(n23531), .ZN(n23530) );
  AND2_X1 U18058 ( .A1(n23526), .A2(net786824), .ZN(n23531) );
  INV_X1 U18059 ( .A(n26018), .ZN(n23526) );
  NAND3_X1 U18060 ( .A1(n23535), .A2(n25588), .A3(n26705), .ZN(n23536) );
  NAND3_X1 U18061 ( .A1(n18193), .A2(n26511), .A3(net720302), .ZN(n23535) );
  INV_X1 U18062 ( .A(n20118), .ZN(net720304) );
  NAND2_X1 U18063 ( .A1(n23538), .A2(n23537), .ZN(n26072) );
  INV_X1 U18064 ( .A(n26209), .ZN(n23537) );
  XNOR2_X1 U18065 ( .A(n26208), .B(net716215), .ZN(n23538) );
  NOR2_X1 U18066 ( .A1(n23539), .A2(net715418), .ZN(n26105) );
  OAI22_X1 U18067 ( .A1(n793), .A2(net715421), .B1(n25282), .B2(net786841), 
        .ZN(n23539) );
  NOR2_X1 U18068 ( .A1(n23540), .A2(n23541), .ZN(n26047) );
  NAND2_X1 U18069 ( .A1(n23542), .A2(n23543), .ZN(n23541) );
  NAND2_X1 U18070 ( .A1(n25420), .A2(net731329), .ZN(n23543) );
  INV_X1 U18071 ( .A(n25946), .ZN(n23542) );
  CLKBUF_X1 U18072 ( .A(net717543), .Z(net755631) );
  OAI21_X1 U18073 ( .B1(n26574), .B2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [12]), .A(n26573), .ZN(n23544) );
  NOR2_X1 U18074 ( .A1(n23545), .A2(n23546), .ZN(n25837) );
  NOR2_X1 U18075 ( .A1(net718134), .A2(n6330), .ZN(n23546) );
  NOR2_X1 U18076 ( .A1(net742037), .A2(n25323), .ZN(n23545) );
  NOR2_X1 U18077 ( .A1(n23547), .A2(net747437), .ZN(net714076) );
  OAI22_X1 U18078 ( .A1(net718337), .A2(n25308), .B1(net718432), .B2(n1718), 
        .ZN(n23547) );
  OAI211_X1 U18079 ( .C1(n22687), .C2(net718133), .A(n23549), .B(n23548), .ZN(
        n25995) );
  OR2_X1 U18080 ( .A1(net765629), .A2(n562), .ZN(n23548) );
  NOR2_X1 U18081 ( .A1(n23550), .A2(n23551), .ZN(n23549) );
  NOR2_X1 U18082 ( .A1(net741958), .A2(n4361), .ZN(n23551) );
  OAI22_X1 U18083 ( .A1(n25354), .A2(net749495), .B1(net765744), .B2(n1742), 
        .ZN(n23550) );
  NOR3_X1 U18084 ( .A1(n25859), .A2(n23552), .A3(n23553), .ZN(n26039) );
  NAND2_X1 U18085 ( .A1(n25856), .A2(n25858), .ZN(n23553) );
  NAND3_X1 U18086 ( .A1(n25857), .A2(net715027), .A3(n25860), .ZN(n23552) );
  NAND3_X1 U18087 ( .A1(n23556), .A2(n23555), .A3(n23554), .ZN(n26096) );
  OR2_X1 U18088 ( .A1(net718337), .A2(n4344), .ZN(n23554) );
  OR2_X1 U18089 ( .A1(net718154), .A2(n1704), .ZN(n23555) );
  AOI22_X1 U18090 ( .A1(net718341), .A2(n24602), .B1(n24275), .B2(n25352), 
        .ZN(n23556) );
  INV_X1 U18091 ( .A(net715180), .ZN(net715175) );
  OAI22_X1 U18092 ( .A1(net767340), .A2(n1678), .B1(net742037), .B2(n5610), 
        .ZN(net715180) );
  NAND2_X1 U18093 ( .A1(n25444), .A2(n23558), .ZN(n25449) );
  INV_X1 U18094 ( .A(n23557), .ZN(n23558) );
  OR2_X1 U18095 ( .A1(n25790), .A2(n24203), .ZN(n23557) );
  NOR2_X1 U18096 ( .A1(n25922), .A2(n23559), .ZN(n25444) );
  NAND2_X1 U18097 ( .A1(n26063), .A2(n24291), .ZN(n23559) );
  NAND3_X1 U18098 ( .A1(n23560), .A2(n23561), .A3(n23562), .ZN(n26113) );
  NAND2_X1 U18099 ( .A1(n24275), .A2(net399701), .ZN(n23562) );
  AOI22_X1 U18100 ( .A1(net715443), .A2(\core_inst/MEMWB_ALUOUT/DFF_5/N3 ), 
        .B1(net755033), .B2(net366478), .ZN(n23560) );
  NAND2_X1 U18101 ( .A1(net718341), .A2(net365826), .ZN(n23561) );
  INV_X1 U18102 ( .A(net712794), .ZN(net712793) );
  INV_X1 U18103 ( .A(n23563), .ZN(n25838) );
  OAI22_X1 U18104 ( .A1(n4400), .A2(n25595), .B1(net717615), .B2(n25324), .ZN(
        n23563) );
  AND2_X1 U18105 ( .A1(net755733), .A2(n23564), .ZN(net733611) );
  NOR2_X1 U18106 ( .A1(n24541), .A2(n24032), .ZN(n23564) );
  NAND2_X1 U18107 ( .A1(n23565), .A2(n23566), .ZN(n26050) );
  OR3_X1 U18108 ( .A1(n25778), .A2(n25777), .A3(net742092), .ZN(n23566) );
  NAND2_X1 U18109 ( .A1(n26144), .A2(net742092), .ZN(n23565) );
  BUF_X1 U18110 ( .A(n23567), .Z(n25578) );
  OAI22_X1 U18111 ( .A1(n26080), .A2(net741686), .B1(net716237), .B2(
        \core_inst/EXMEM_NPC/DFF_27/N3 ), .ZN(n23567) );
  NOR2_X1 U18112 ( .A1(n26000), .A2(net714382), .ZN(net714502) );
  OAI21_X1 U18113 ( .B1(n25996), .B2(net749977), .A(n23568), .ZN(net714501) );
  AOI22_X1 U18114 ( .A1(n26226), .A2(net767234), .B1(n26224), .B2(n26136), 
        .ZN(n23568) );
  NAND3_X1 U18115 ( .A1(n23569), .A2(n23570), .A3(n23571), .ZN(n26080) );
  NAND2_X1 U18116 ( .A1(n25390), .A2(n14769), .ZN(n23571) );
  NAND2_X1 U18117 ( .A1(net718340), .A2(n24783), .ZN(n23570) );
  AOI22_X1 U18118 ( .A1(net715443), .A2(\core_inst/MEMWB_ALUOUT/DFF_27/N3 ), 
        .B1(net715445), .B2(n561), .ZN(n23569) );
  NOR2_X1 U18119 ( .A1(n23573), .A2(n23572), .ZN(n26144) );
  OAI22_X1 U18120 ( .A1(n25787), .A2(net717570), .B1(n26071), .B2(n25782), 
        .ZN(n23572) );
  OAI22_X1 U18121 ( .A1(net713633), .A2(n25781), .B1(n23574), .B2(net755207), 
        .ZN(n23573) );
  NAND2_X1 U18122 ( .A1(n25578), .A2(net717570), .ZN(n23574) );
  XNOR2_X1 U18123 ( .A(n23575), .B(net716223), .ZN(n23576) );
  NAND2_X1 U18124 ( .A1(n25827), .A2(n25826), .ZN(n23575) );
  INV_X1 U18125 ( .A(n23577), .ZN(n25576) );
  MUX2_X1 U18126 ( .A(n26112), .B(\core_inst/EXMEM_NPC/DFF_6/N3 ), .S(
        net741686), .Z(n23577) );
  NAND2_X1 U18127 ( .A1(n26027), .A2(n24558), .ZN(net763705) );
  OAI222_X1 U18128 ( .A1(net780556), .A2(n24555), .B1(n24402), .B2(net714494), 
        .C1(net713633), .C2(n24276), .ZN(n25378) );
  NAND3_X1 U18129 ( .A1(n23578), .A2(n23579), .A3(n23580), .ZN(n26112) );
  NAND2_X1 U18130 ( .A1(n25390), .A2(n25342), .ZN(n23580) );
  NAND2_X1 U18131 ( .A1(net718341), .A2(n24780), .ZN(n23579) );
  AOI22_X1 U18132 ( .A1(net715443), .A2(\core_inst/MEMWB_ALUOUT/DFF_6/N3 ), 
        .B1(net715445), .B2(n5729), .ZN(n23578) );
  AOI211_X2 U18133 ( .C1(n26195), .C2(n26251), .A(n23581), .B(n23582), .ZN(
        n26250) );
  NOR3_X1 U18134 ( .A1(n23583), .A2(n26194), .A3(n24301), .ZN(n23582) );
  INV_X1 U18135 ( .A(n26192), .ZN(n23583) );
  INV_X1 U18136 ( .A(n26191), .ZN(n23581) );
  NAND4_X1 U18137 ( .A1(n23584), .A2(n23585), .A3(n23586), .A4(n23587), .ZN(
        n25749) );
  XOR2_X1 U18138 ( .A(net366410), .B(n1651), .Z(n23587) );
  XOR2_X1 U18139 ( .A(net342954), .B(n5174), .Z(n23586) );
  XOR2_X1 U18140 ( .A(n25590), .B(n5598), .Z(n23585) );
  NOR2_X1 U18141 ( .A1(n23588), .A2(n23589), .ZN(n23584) );
  XNOR2_X1 U18142 ( .A(net366411), .B(n5613), .ZN(n23589) );
  XOR2_X1 U18143 ( .A(net342961), .B(n18053), .Z(n23588) );
  NAND4_X1 U18144 ( .A1(n23590), .A2(n23591), .A3(net716231), .A4(n25756), 
        .ZN(n25757) );
  INV_X1 U18145 ( .A(n23594), .ZN(n23591) );
  CLKBUF_X1 U18146 ( .A(n25755), .Z(n23594) );
  NOR2_X1 U18147 ( .A1(n23592), .A2(n23593), .ZN(n23590) );
  INV_X1 U18148 ( .A(n25754), .ZN(n23593) );
  INV_X1 U18149 ( .A(n25753), .ZN(n23592) );
  MUX2_X1 U18150 ( .A(n23595), .B(n26023), .S(net717510), .Z(net713977) );
  OR2_X1 U18151 ( .A1(n25778), .A2(n25777), .ZN(n23595) );
  NOR2_X1 U18152 ( .A1(n23596), .A2(n23597), .ZN(n25853) );
  NOR2_X1 U18153 ( .A1(net741959), .A2(n4382), .ZN(n23597) );
  OAI22_X1 U18154 ( .A1(net749972), .A2(n1702), .B1(net767205), .B2(n25309), 
        .ZN(n23596) );
  NAND3_X1 U18155 ( .A1(net736610), .A2(n23598), .A3(net736609), .ZN(n26108)
         );
  CLKBUF_X1 U18156 ( .A(net718341), .Z(net750031) );
  NAND2_X1 U18157 ( .A1(n25390), .A2(n17664), .ZN(n23598) );
  OR2_X1 U18158 ( .A1(n23599), .A2(n25379), .ZN(n23979) );
  NOR2_X1 U18159 ( .A1(n25823), .A2(net755228), .ZN(n23599) );
  INV_X1 U18160 ( .A(net742146), .ZN(net755228) );
  NOR2_X1 U18161 ( .A1(n23600), .A2(n23601), .ZN(n25836) );
  AND2_X1 U18162 ( .A1(n24320), .A2(n25327), .ZN(n23601) );
  OAI22_X1 U18163 ( .A1(n1732), .A2(net717106), .B1(net749495), .B2(n4404), 
        .ZN(n23600) );
  XNOR2_X1 U18164 ( .A(n23602), .B(net716215), .ZN(n24028) );
  NAND3_X1 U18165 ( .A1(n23326), .A2(n26048), .A3(n26049), .ZN(n23602) );
  INV_X1 U18166 ( .A(net713966), .ZN(net714542) );
  XNOR2_X1 U18167 ( .A(n26034), .B(n23603), .ZN(n24382) );
  NOR2_X1 U18168 ( .A1(n24324), .A2(n24176), .ZN(n23603) );
  NOR2_X1 U18169 ( .A1(n23604), .A2(n24192), .ZN(n25937) );
  XNOR2_X1 U18170 ( .A(net742241), .B(net716215), .ZN(n23604) );
  NAND3_X1 U18171 ( .A1(n23605), .A2(n23606), .A3(n23607), .ZN(n26195) );
  NAND3_X1 U18172 ( .A1(net713692), .A2(net742324), .A3(n23610), .ZN(n23607)
         );
  INV_X1 U18173 ( .A(n24285), .ZN(n23610) );
  NAND2_X1 U18174 ( .A1(net749306), .A2(n24091), .ZN(n23606) );
  NAND3_X1 U18175 ( .A1(n23608), .A2(n23609), .A3(net713692), .ZN(n23605) );
  NOR2_X1 U18176 ( .A1(n26182), .A2(n26183), .ZN(n23609) );
  OAI22_X1 U18177 ( .A1(n24170), .A2(net749832), .B1(net713711), .B2(net755090), .ZN(n23608) );
  OR2_X1 U18178 ( .A1(n24273), .A2(n23611), .ZN(n25502) );
  OAI21_X1 U18179 ( .B1(n23612), .B2(n23614), .A(n24557), .ZN(n23611) );
  AOI21_X1 U18180 ( .B1(net714947), .B2(net728158), .A(net714724), .ZN(n23614)
         );
  NAND2_X1 U18181 ( .A1(n23613), .A2(n23023), .ZN(n23612) );
  NOR2_X1 U18182 ( .A1(n24353), .A2(n26118), .ZN(n23613) );
  NAND2_X1 U18183 ( .A1(n24193), .A2(n25337), .ZN(n23615) );
  OAI22_X1 U18184 ( .A1(net780584), .A2(net740655), .B1(net717106), .B2(n1720), 
        .ZN(n23616) );
  OAI22_X1 U18185 ( .A1(net767341), .A2(n23271), .B1(net717615), .B2(n5595), 
        .ZN(n23617) );
  NOR2_X1 U18186 ( .A1(n23616), .A2(n23617), .ZN(n23618) );
  NAND2_X1 U18187 ( .A1(n23615), .A2(n23618), .ZN(net713561) );
  INV_X1 U18188 ( .A(n23619), .ZN(n25844) );
  OAI22_X1 U18189 ( .A1(n1659), .A2(net767340), .B1(net742037), .B2(n5186), 
        .ZN(n23619) );
  NOR2_X1 U18190 ( .A1(n23620), .A2(net768639), .ZN(n25392) );
  OAI22_X1 U18191 ( .A1(net742209), .A2(n25359), .B1(net717718), .B2(n24609), 
        .ZN(n23620) );
  NOR2_X1 U18192 ( .A1(n23621), .A2(n23622), .ZN(net724632) );
  NOR2_X1 U18193 ( .A1(net750086), .A2(n4364), .ZN(n23622) );
  OAI22_X1 U18194 ( .A1(net767205), .A2(n25350), .B1(net749972), .B2(n1728), 
        .ZN(n23621) );
  NAND2_X1 U18195 ( .A1(n23623), .A2(net769389), .ZN(net715656) );
  INV_X1 U18196 ( .A(net718033), .ZN(net769389) );
  NAND2_X1 U18197 ( .A1(net740075), .A2(net715666), .ZN(n23623) );
  NAND2_X1 U18198 ( .A1(n26532), .A2(n23624), .ZN(n25922) );
  NOR2_X1 U18199 ( .A1(n26531), .A2(n26062), .ZN(n23624) );
  OAI22_X1 U18200 ( .A1(n24543), .A2(n24572), .B1(net713151), .B2(net755013), 
        .ZN(n25792) );
  CLKBUF_X1 U18201 ( .A(net717543), .Z(net755013) );
  NAND2_X1 U18202 ( .A1(n23625), .A2(net714873), .ZN(n25377) );
  AOI22_X1 U18203 ( .A1(net750025), .A2(net713773), .B1(net749500), .B2(
        net718391), .ZN(n23625) );
  XNOR2_X1 U18204 ( .A(net366411), .B(net749230), .ZN(net715784) );
  XNOR2_X1 U18205 ( .A(net342963), .B(net749551), .ZN(net715783) );
  OAI222_X1 U18206 ( .A1(net749926), .A2(n5611), .B1(net714943), .B2(n4410), 
        .C1(net765744), .C2(n1744), .ZN(n23626) );
  NAND2_X1 U18207 ( .A1(n24320), .A2(net740710), .ZN(n23627) );
  OAI21_X1 U18208 ( .B1(net718134), .B2(net89402), .A(n23627), .ZN(n23628) );
  OR2_X1 U18209 ( .A1(n23626), .A2(n23628), .ZN(n25887) );
  NAND2_X1 U18210 ( .A1(n25587), .A2(n24576), .ZN(net715050) );
  NAND4_X1 U18211 ( .A1(n23629), .A2(n23630), .A3(n23631), .A4(n23632), .ZN(
        n25987) );
  NAND3_X1 U18212 ( .A1(net749260), .A2(net749534), .A3(n22673), .ZN(n23632)
         );
  NAND2_X1 U18213 ( .A1(net717875), .A2(n25786), .ZN(n23631) );
  NAND2_X1 U18214 ( .A1(n24341), .A2(n25785), .ZN(n23630) );
  NAND2_X1 U18215 ( .A1(net755240), .A2(n24190), .ZN(n23629) );
  NAND2_X1 U18216 ( .A1(n23633), .A2(n23634), .ZN(n25832) );
  NOR2_X1 U18217 ( .A1(n23635), .A2(n23637), .ZN(n23634) );
  AND2_X1 U18218 ( .A1(net749274), .A2(n25318), .ZN(n23637) );
  OAI22_X1 U18219 ( .A1(net717106), .A2(n1724), .B1(net780584), .B2(n25311), 
        .ZN(n23635) );
  INV_X1 U18220 ( .A(n23636), .ZN(n23633) );
  OAI22_X1 U18221 ( .A1(n23264), .A2(net767341), .B1(net715058), .B2(n756), 
        .ZN(n23636) );
  NAND3_X1 U18222 ( .A1(n25772), .A2(n23638), .A3(n25774), .ZN(n26040) );
  AND2_X1 U18223 ( .A1(n25771), .A2(n25770), .ZN(n23638) );
  NOR2_X1 U18224 ( .A1(n23639), .A2(n23640), .ZN(n25772) );
  OAI22_X1 U18225 ( .A1(net762729), .A2(net746701), .B1(net713151), .B2(n25789), .ZN(n23640) );
  OAI22_X1 U18226 ( .A1(net750090), .A2(net714871), .B1(n24276), .B2(net713707), .ZN(n23639) );
  NAND4_X1 U18227 ( .A1(n23641), .A2(n25940), .A3(net715050), .A4(n25935), 
        .ZN(n25846) );
  NAND2_X1 U18228 ( .A1(n24197), .A2(n26041), .ZN(n23641) );
  NAND2_X1 U18229 ( .A1(n25420), .A2(net731327), .ZN(n23642) );
  NAND2_X2 U18230 ( .A1(n23643), .A2(n23644), .ZN(net713607) );
  OR2_X1 U18231 ( .A1(net787528), .A2(n6740), .ZN(n23644) );
  NAND2_X1 U18232 ( .A1(n26086), .A2(net787512), .ZN(n23643) );
  NAND3_X1 U18233 ( .A1(net715536), .A2(n23645), .A3(n23646), .ZN(n26086) );
  NAND2_X1 U18234 ( .A1(n25390), .A2(n25340), .ZN(n23646) );
  NAND2_X1 U18235 ( .A1(net718341), .A2(n25337), .ZN(n23645) );
  CLKBUF_X1 U18236 ( .A(net715445), .Z(net750111) );
  NAND2_X1 U18237 ( .A1(n25940), .A2(n23647), .ZN(n26067) );
  NAND2_X1 U18238 ( .A1(n24031), .A2(n25936), .ZN(n23647) );
  AND3_X1 U18239 ( .A1(n25776), .A2(n23648), .A3(n25775), .ZN(n24545) );
  AND2_X1 U18240 ( .A1(n25773), .A2(n25774), .ZN(n23648) );
  OAI21_X1 U18241 ( .B1(n26132), .B2(n24290), .A(n23649), .ZN(n25382) );
  AOI21_X1 U18242 ( .B1(n25379), .B2(n23650), .A(n24538), .ZN(n23649) );
  AOI21_X1 U18243 ( .B1(n25898), .B2(n23977), .A(n24202), .ZN(n23650) );
  NOR2_X1 U18244 ( .A1(n23651), .A2(net715586), .ZN(n26184) );
  OAI22_X1 U18245 ( .A1(n4343), .A2(n25595), .B1(n24815), .B2(net738474), .ZN(
        n23651) );
  XNOR2_X1 U18246 ( .A(n23652), .B(n26509), .ZN(net712976) );
  OAI21_X1 U18247 ( .B1(n23653), .B2(n24542), .A(n23654), .ZN(n23652) );
  AOI21_X1 U18248 ( .B1(n24563), .B2(n26247), .A(n26238), .ZN(n23654) );
  NAND3_X1 U18249 ( .A1(n23655), .A2(n26248), .A3(n25504), .ZN(n23653) );
  NAND3_X1 U18250 ( .A1(n23656), .A2(n22830), .A3(n26250), .ZN(n23655) );
  NAND3_X1 U18251 ( .A1(n26236), .A2(n23657), .A3(n26237), .ZN(n23656) );
  AND2_X1 U18252 ( .A1(n26251), .A2(n24843), .ZN(n23657) );
  NOR2_X1 U18253 ( .A1(n24548), .A2(n23966), .ZN(n23658) );
  NAND2_X1 U18254 ( .A1(n23659), .A2(n26250), .ZN(n26248) );
  NOR4_X1 U18255 ( .A1(n26220), .A2(n23660), .A3(n23661), .A4(n23662), .ZN(
        n23659) );
  NAND2_X1 U18256 ( .A1(n26219), .A2(n26218), .ZN(n23662) );
  NAND3_X1 U18257 ( .A1(n26217), .A2(n26216), .A3(n26215), .ZN(n23661) );
  INV_X1 U18258 ( .A(n26253), .ZN(n23660) );
  NAND2_X1 U18259 ( .A1(n23663), .A2(n23664), .ZN(n25765) );
  NAND3_X1 U18260 ( .A1(n25772), .A2(n23665), .A3(n25774), .ZN(n23664) );
  AND3_X1 U18261 ( .A1(n25771), .A2(net714275), .A3(n25770), .ZN(n23665) );
  NAND3_X1 U18262 ( .A1(n24331), .A2(n25371), .A3(net714309), .ZN(n23663) );
  INV_X1 U18263 ( .A(n23666), .ZN(n24374) );
  OAI22_X1 U18264 ( .A1(n23265), .A2(net767340), .B1(net749972), .B2(n1698), 
        .ZN(n23666) );
  NOR2_X1 U18265 ( .A1(n23668), .A2(n23669), .ZN(net729292) );
  NOR2_X1 U18266 ( .A1(n26076), .A2(net713728), .ZN(n23669) );
  AND2_X1 U18267 ( .A1(n26076), .A2(net767168), .ZN(n23668) );
  NAND3_X1 U18268 ( .A1(n23667), .A2(net717091), .A3(n26075), .ZN(net729291)
         );
  NAND2_X1 U18269 ( .A1(net713813), .A2(n26073), .ZN(n23667) );
  NOR2_X1 U18270 ( .A1(net715695), .A2(net749843), .ZN(net715668) );
  AND2_X1 U18271 ( .A1(n23670), .A2(n23671), .ZN(net737707) );
  NAND3_X1 U18272 ( .A1(n23680), .A2(n23681), .A3(n23679), .ZN(n23671) );
  NOR2_X1 U18273 ( .A1(n24568), .A2(n23688), .ZN(n23681) );
  NOR3_X1 U18274 ( .A1(n23676), .A2(n23677), .A3(n23678), .ZN(n23670) );
  OAI211_X1 U18275 ( .C1(n23672), .C2(n23673), .A(n23675), .B(n23674), .ZN(
        net714140) );
  AOI21_X1 U18276 ( .B1(n23678), .B2(n23677), .A(net713154), .ZN(n23674) );
  NOR2_X1 U18277 ( .A1(n22837), .A2(n23685), .ZN(n23678) );
  NAND2_X1 U18278 ( .A1(n24317), .A2(n24138), .ZN(n23685) );
  NAND2_X1 U18279 ( .A1(n23676), .A2(n23677), .ZN(n23675) );
  AOI211_X1 U18280 ( .C1(net714164), .C2(n23684), .A(n23688), .B(n23682), .ZN(
        n23676) );
  NOR2_X1 U18281 ( .A1(n24278), .A2(n24305), .ZN(n23688) );
  AND2_X1 U18282 ( .A1(n26067), .A2(n23686), .ZN(n23684) );
  NAND4_X1 U18283 ( .A1(n23679), .A2(net742326), .A3(n24138), .A4(n23677), 
        .ZN(n23673) );
  XNOR2_X1 U18284 ( .A(n23683), .B(n24033), .ZN(n23677) );
  INV_X1 U18285 ( .A(n23952), .ZN(n23683) );
  INV_X1 U18286 ( .A(n22837), .ZN(n23679) );
  NOR2_X1 U18287 ( .A1(n23687), .A2(n24549), .ZN(n23682) );
  NAND2_X1 U18288 ( .A1(n26067), .A2(n23686), .ZN(n23687) );
  OR2_X1 U18289 ( .A1(n24265), .A2(n24029), .ZN(n23686) );
  INV_X1 U18290 ( .A(n23680), .ZN(n23672) );
  NOR2_X1 U18291 ( .A1(n26069), .A2(net714157), .ZN(n23680) );
  NOR2_X1 U18292 ( .A1(n23689), .A2(n23690), .ZN(n25403) );
  NOR2_X1 U18293 ( .A1(n24033), .A2(n24276), .ZN(n23690) );
  NAND3_X1 U18294 ( .A1(n25884), .A2(n23691), .A3(n23692), .ZN(n23689) );
  OR2_X1 U18295 ( .A1(n25600), .A2(net749685), .ZN(n23692) );
  NAND2_X1 U18296 ( .A1(net749489), .A2(n24577), .ZN(n23691) );
  MUX2_X1 U18297 ( .A(net715706), .B(net715707), .S(s_MEMWB_IR[27]), .Z(
        net715834) );
  AOI21_X1 U18298 ( .B1(n23693), .B2(n25981), .A(n25941), .ZN(net712882) );
  NOR2_X1 U18299 ( .A1(n24571), .A2(net750238), .ZN(n23693) );
  NOR2_X1 U18300 ( .A1(n23694), .A2(n23695), .ZN(n26088) );
  OAI22_X1 U18301 ( .A1(net715420), .A2(n25307), .B1(net742413), .B2(n1698), 
        .ZN(n23695) );
  OAI22_X1 U18302 ( .A1(net715422), .A2(n4379), .B1(n716), .B2(net715421), 
        .ZN(n23694) );
  NAND2_X1 U18303 ( .A1(n23696), .A2(n23697), .ZN(n25369) );
  OR2_X1 U18304 ( .A1(n25370), .A2(n25746), .ZN(n23697) );
  XNOR2_X1 U18305 ( .A(net718081), .B(s_MEMWB_IR[19]), .ZN(n23696) );
  NOR2_X1 U18306 ( .A1(n23698), .A2(n23699), .ZN(n24259) );
  OAI22_X1 U18307 ( .A1(net762729), .A2(net713607), .B1(n25789), .B2(net713564), .ZN(n23699) );
  OAI22_X1 U18308 ( .A1(n26193), .A2(net749902), .B1(net780556), .B2(net750032), .ZN(n23698) );
  INV_X1 U18309 ( .A(n23700), .ZN(n24397) );
  OAI22_X1 U18310 ( .A1(n24342), .A2(net767209), .B1(n23701), .B2(net713154), 
        .ZN(n23700) );
  XNOR2_X1 U18311 ( .A(n25447), .B(n23702), .ZN(n23701) );
  AND2_X1 U18312 ( .A1(n24308), .A2(n26036), .ZN(n23702) );
  AOI222_X1 U18313 ( .A1(net714249), .A2(net767206), .B1(n26148), .B2(n24341), 
        .C1(n23969), .C2(net750057), .ZN(n25425) );
  NAND2_X1 U18314 ( .A1(net729186), .A2(n25413), .ZN(net729185) );
  NAND2_X1 U18315 ( .A1(n23704), .A2(n24566), .ZN(net729177) );
  NOR2_X1 U18316 ( .A1(n23705), .A2(n23706), .ZN(n23704) );
  NAND2_X1 U18317 ( .A1(n23709), .A2(n23710), .ZN(n23706) );
  OR2_X1 U18318 ( .A1(n24328), .A2(net749709), .ZN(n23710) );
  OR2_X1 U18319 ( .A1(net767209), .A2(n23703), .ZN(n23709) );
  NAND2_X1 U18320 ( .A1(n25900), .A2(n25899), .ZN(n23703) );
  OAI222_X1 U18321 ( .A1(n24330), .A2(net714267), .B1(n26046), .B2(net713897), 
        .C1(n23707), .C2(n23708), .ZN(n23705) );
  NAND2_X1 U18322 ( .A1(n26045), .A2(n26044), .ZN(n23708) );
  NOR2_X1 U18323 ( .A1(n23712), .A2(n23711), .ZN(n26089) );
  OAI22_X1 U18324 ( .A1(n5187), .A2(net742209), .B1(n4382), .B2(net717719), 
        .ZN(n23711) );
  OAI22_X1 U18325 ( .A1(n1702), .A2(net715419), .B1(net742223), .B2(n25309), 
        .ZN(n23712) );
  MUX2_X2 U18326 ( .A(n23713), .B(n23714), .S(net742092), .Z(net713870) );
  INV_X1 U18327 ( .A(n25998), .ZN(n23714) );
  NAND4_X1 U18328 ( .A1(n23715), .A2(net715333), .A3(n23716), .A4(n23717), 
        .ZN(n25998) );
  NAND2_X1 U18329 ( .A1(net713701), .A2(n25786), .ZN(n23717) );
  NAND2_X1 U18330 ( .A1(net713905), .A2(n24190), .ZN(n23716) );
  NAND2_X1 U18331 ( .A1(n24345), .A2(n25785), .ZN(n23715) );
  NOR2_X1 U18332 ( .A1(n25600), .A2(net742473), .ZN(net717780) );
  NOR2_X1 U18333 ( .A1(n24267), .A2(n24525), .ZN(net717779) );
  NOR2_X1 U18334 ( .A1(net750203), .A2(n24548), .ZN(net717778) );
  NAND3_X1 U18335 ( .A1(n23718), .A2(n23719), .A3(n23720), .ZN(n25997) );
  NAND2_X1 U18336 ( .A1(n25909), .A2(n24206), .ZN(n23720) );
  NAND2_X1 U18337 ( .A1(net713672), .A2(net750255), .ZN(n23719) );
  AOI21_X1 U18338 ( .B1(net749454), .B2(n25788), .A(n25815), .ZN(n23718) );
  OR2_X1 U18339 ( .A1(net742413), .A2(n1732), .ZN(n23721) );
  AOI22_X1 U18340 ( .A1(net718341), .A2(n25327), .B1(n24275), .B2(n11928), 
        .ZN(n23722) );
  OAI211_X1 U18341 ( .C1(net715420), .C2(n4404), .A(n23721), .B(n23722), .ZN(
        n26091) );
  INV_X1 U18342 ( .A(n23723), .ZN(n25822) );
  XNOR2_X1 U18343 ( .A(n23724), .B(net716215), .ZN(n26035) );
  NAND2_X1 U18344 ( .A1(n25822), .A2(n23725), .ZN(n23724) );
  NOR2_X1 U18345 ( .A1(net715221), .A2(n25821), .ZN(n23725) );
  NOR2_X1 U18346 ( .A1(n23726), .A2(n25505), .ZN(n26150) );
  NAND3_X1 U18347 ( .A1(n23822), .A2(n23727), .A3(n25416), .ZN(n23726) );
  NAND3_X1 U18348 ( .A1(n25752), .A2(net786837), .A3(net725586), .ZN(n23727)
         );
  NAND2_X1 U18349 ( .A1(net749922), .A2(net740639), .ZN(n25509) );
  NAND2_X1 U18350 ( .A1(n23730), .A2(n25760), .ZN(net715586) );
  AND2_X1 U18351 ( .A1(net715524), .A2(n23728), .ZN(n23730) );
  NAND3_X1 U18352 ( .A1(n23729), .A2(net742282), .A3(net715591), .ZN(n23728)
         );
  NOR2_X1 U18353 ( .A1(net715592), .A2(net750079), .ZN(n23729) );
  NAND3_X1 U18354 ( .A1(n23731), .A2(n23732), .A3(n23733), .ZN(n25471) );
  NOR2_X1 U18355 ( .A1(n26061), .A2(n24322), .ZN(n23733) );
  NOR3_X1 U18356 ( .A1(n24300), .A2(n26172), .A3(n24321), .ZN(n23731) );
  NAND2_X1 U18357 ( .A1(n23735), .A2(net732762), .ZN(n26406) );
  NAND3_X1 U18358 ( .A1(n23734), .A2(n23736), .A3(net717074), .ZN(n23735) );
  AND3_X1 U18359 ( .A1(n23737), .A2(n24310), .A3(net748264), .ZN(n23736) );
  INV_X1 U18360 ( .A(net712468), .ZN(net748264) );
  AND2_X1 U18361 ( .A1(net750287), .A2(net728314), .ZN(n23737) );
  NOR2_X1 U18362 ( .A1(n24425), .A2(n25471), .ZN(n23734) );
  NAND2_X1 U18363 ( .A1(n26075), .A2(n23738), .ZN(net713448) );
  NOR3_X1 U18364 ( .A1(n23739), .A2(n23740), .A3(n23741), .ZN(n23738) );
  AND3_X1 U18365 ( .A1(net717547), .A2(net749428), .A3(n26209), .ZN(n23741) );
  INV_X1 U18366 ( .A(n25943), .ZN(n23740) );
  NOR3_X1 U18367 ( .A1(net714113), .A2(net749945), .A3(n24525), .ZN(n23739) );
  NAND2_X1 U18368 ( .A1(n25749), .A2(n23742), .ZN(n24262) );
  NOR3_X1 U18369 ( .A1(n23743), .A2(n23744), .A3(n23745), .ZN(n23742) );
  NAND3_X1 U18370 ( .A1(n23746), .A2(n23747), .A3(n23748), .ZN(n23745) );
  XNOR2_X1 U18371 ( .A(n1665), .B(n5598), .ZN(n23748) );
  XNOR2_X1 U18372 ( .A(n1668), .B(n1651), .ZN(n23747) );
  XNOR2_X1 U18373 ( .A(n1666), .B(n5174), .ZN(n23746) );
  XNOR2_X1 U18374 ( .A(net342852), .B(n5613), .ZN(n23744) );
  XOR2_X1 U18375 ( .A(net342960), .B(n18053), .Z(n23743) );
  XNOR2_X1 U18376 ( .A(net718069), .B(n25582), .ZN(n23749) );
  XNOR2_X1 U18377 ( .A(n25592), .B(n25593), .ZN(n23750) );
  XOR2_X1 U18378 ( .A(net718070), .B(s_MEMWB_IR[18]), .Z(n23751) );
  NAND3_X1 U18379 ( .A1(n23752), .A2(n23753), .A3(n23754), .ZN(n26111) );
  NAND2_X1 U18380 ( .A1(net750135), .A2(\core_inst/MEMWB_ALUOUT/DFF_10/N3 ), 
        .ZN(n23754) );
  OAI21_X1 U18381 ( .B1(n23755), .B2(n23756), .A(net796122), .ZN(n23753) );
  NOR2_X1 U18382 ( .A1(n4415), .A2(net749369), .ZN(n23756) );
  NOR2_X1 U18383 ( .A1(net749951), .A2(n4416), .ZN(n23755) );
  NAND2_X1 U18384 ( .A1(n25390), .A2(n17665), .ZN(n23752) );
  OAI22_X1 U18385 ( .A1(n23758), .A2(n25974), .B1(n24530), .B2(n23759), .ZN(
        net728481) );
  NOR2_X1 U18386 ( .A1(n23757), .A2(n23760), .ZN(n23759) );
  NAND2_X1 U18387 ( .A1(n23761), .A2(net714006), .ZN(n23760) );
  NOR3_X1 U18388 ( .A1(n24319), .A2(n24089), .A3(n23023), .ZN(n23761) );
  NOR2_X1 U18389 ( .A1(net720121), .A2(n25372), .ZN(n23757) );
  NAND2_X1 U18390 ( .A1(n23762), .A2(n26256), .ZN(n23758) );
  NOR2_X1 U18391 ( .A1(n25405), .A2(n25874), .ZN(n23762) );
  NAND2_X1 U18392 ( .A1(n24031), .A2(n25936), .ZN(n23764) );
  AND2_X1 U18393 ( .A1(n24350), .A2(n23765), .ZN(n23763) );
  OR2_X1 U18394 ( .A1(n23952), .A2(n24033), .ZN(n23765) );
  NOR2_X1 U18395 ( .A1(net715015), .A2(n23766), .ZN(n24561) );
  NAND3_X1 U18396 ( .A1(n23767), .A2(net718024), .A3(n26219), .ZN(n25985) );
  INV_X1 U18397 ( .A(net755260), .ZN(net718024) );
  AOI22_X1 U18398 ( .A1(net750238), .A2(n25788), .B1(net713753), .B2(n22673), 
        .ZN(n23767) );
  AND2_X1 U18399 ( .A1(net713845), .A2(\core_inst/MEMWB_ALUOUT/DFF_11/N3 ), 
        .ZN(n23769) );
  OAI22_X1 U18400 ( .A1(net749926), .A2(n25325), .B1(net718361), .B2(n17859), 
        .ZN(n23768) );
  XNOR2_X1 U18401 ( .A(n23770), .B(net741307), .ZN(n25587) );
  NAND2_X1 U18402 ( .A1(n25844), .A2(n25843), .ZN(n23770) );
  NAND3_X1 U18403 ( .A1(n1668), .A2(n1666), .A3(n1665), .ZN(n23771) );
  NAND2_X1 U18404 ( .A1(n25861), .A2(n23772), .ZN(n25758) );
  MUX2_X1 U18405 ( .A(n26098), .B(\core_inst/EXMEM_NPC/DFF_0/N3 ), .S(
        net741686), .Z(n23772) );
  NAND3_X1 U18406 ( .A1(n23773), .A2(n25758), .A3(n25757), .ZN(n24314) );
  XNOR2_X1 U18407 ( .A(n26150), .B(net716215), .ZN(n23773) );
  NAND2_X1 U18408 ( .A1(n23775), .A2(n23776), .ZN(n26098) );
  AOI22_X1 U18409 ( .A1(n23774), .A2(\core_inst/MEMWB_ALUOUT/DFF_0/N3 ), .B1(
        n23777), .B2(net715460), .ZN(n23776) );
  NOR2_X1 U18410 ( .A1(net749951), .A2(n4422), .ZN(n23777) );
  NOR2_X1 U18411 ( .A1(net749664), .A2(net715460), .ZN(n23774) );
  AOI21_X1 U18412 ( .B1(net718341), .B2(n24781), .A(n23778), .ZN(n23775) );
  NOR3_X1 U18413 ( .A1(net715460), .A2(net749369), .A3(n1537), .ZN(n23778) );
  NAND3_X1 U18414 ( .A1(n23781), .A2(n23782), .A3(n23783), .ZN(n23780) );
  NAND2_X1 U18415 ( .A1(n26018), .A2(n23788), .ZN(n23783) );
  INV_X1 U18416 ( .A(n24339), .ZN(n23788) );
  AOI21_X1 U18417 ( .B1(n23784), .B2(n24538), .A(n23785), .ZN(n23782) );
  NAND3_X1 U18418 ( .A1(net749720), .A2(n24348), .A3(n23784), .ZN(n23781) );
  NOR2_X1 U18419 ( .A1(n25934), .A2(net755086), .ZN(n23784) );
  INV_X1 U18420 ( .A(n22844), .ZN(net749720) );
  OAI21_X1 U18421 ( .B1(net738840), .B2(n24568), .A(n23786), .ZN(n23779) );
  NOR2_X1 U18422 ( .A1(n23787), .A2(n24339), .ZN(n23786) );
  INV_X1 U18423 ( .A(n23785), .ZN(n23787) );
  XNOR2_X1 U18424 ( .A(n23789), .B(n24548), .ZN(n23785) );
  XOR2_X1 U18425 ( .A(n25903), .B(net716215), .Z(n23789) );
  XOR2_X1 U18426 ( .A(n25586), .B(n24356), .Z(net745684) );
  NAND2_X1 U18427 ( .A1(n23794), .A2(n23795), .ZN(net745672) );
  NAND2_X1 U18428 ( .A1(n23796), .A2(net714016), .ZN(n23795) );
  OAI21_X1 U18429 ( .B1(n23797), .B2(net734346), .A(n23790), .ZN(n23796) );
  NOR2_X1 U18430 ( .A1(n23798), .A2(net728159), .ZN(n23797) );
  AND2_X1 U18431 ( .A1(n24086), .A2(net728158), .ZN(n23798) );
  NAND3_X1 U18432 ( .A1(net713467), .A2(n23799), .A3(net745679), .ZN(n23794)
         );
  INV_X1 U18433 ( .A(net714016), .ZN(net745681) );
  NAND2_X1 U18434 ( .A1(n23791), .A2(n23790), .ZN(net714016) );
  INV_X1 U18435 ( .A(n24200), .ZN(n23790) );
  NAND3_X1 U18436 ( .A1(n23792), .A2(n23793), .A3(n24349), .ZN(n23791) );
  INV_X1 U18437 ( .A(n26118), .ZN(n23793) );
  INV_X1 U18438 ( .A(n24353), .ZN(n23792) );
  OR2_X1 U18439 ( .A1(n25438), .A2(net728159), .ZN(n23799) );
  NOR2_X1 U18440 ( .A1(n25405), .A2(n25874), .ZN(net713469) );
  NAND3_X1 U18441 ( .A1(n24529), .A2(net714006), .A3(n25365), .ZN(net714337)
         );
  NOR2_X1 U18442 ( .A1(net720121), .A2(n25372), .ZN(net755783) );
  NAND3_X1 U18443 ( .A1(n23801), .A2(n23802), .A3(n23800), .ZN(n26084) );
  NAND2_X1 U18444 ( .A1(net718341), .A2(n24605), .ZN(n23800) );
  NAND2_X1 U18445 ( .A1(n25390), .A2(n25341), .ZN(n23802) );
  AOI22_X1 U18446 ( .A1(net749408), .A2(n600), .B1(net715443), .B2(
        \core_inst/MEMWB_ALUOUT/DFF_26/N3 ), .ZN(n23801) );
  NAND3_X1 U18447 ( .A1(n24374), .A2(n23803), .A3(n23804), .ZN(n26204) );
  INV_X1 U18448 ( .A(n24376), .ZN(n23804) );
  INV_X1 U18449 ( .A(n24375), .ZN(n23803) );
  AND2_X2 U18450 ( .A1(n23970), .A2(n23805), .ZN(n24541) );
  XNOR2_X1 U18451 ( .A(n26204), .B(net716221), .ZN(n23805) );
  NAND3_X1 U18452 ( .A1(n23806), .A2(n23807), .A3(n25787), .ZN(n26023) );
  NAND2_X1 U18453 ( .A1(net749306), .A2(n22673), .ZN(n23807) );
  AOI21_X1 U18454 ( .B1(net749343), .B2(n25788), .A(n25815), .ZN(n23806) );
  OR3_X1 U18455 ( .A1(n23811), .A2(net714122), .A3(n23808), .ZN(net745868) );
  AOI21_X1 U18456 ( .B1(net740526), .B2(n23809), .A(n23812), .ZN(n23811) );
  OAI21_X1 U18457 ( .B1(n23811), .B2(net714122), .A(n23808), .ZN(net745867) );
  XNOR2_X1 U18458 ( .A(n26071), .B(net742492), .ZN(n23808) );
  CLKBUF_X1 U18459 ( .A(net749636), .Z(net742492) );
  NAND2_X1 U18460 ( .A1(n23810), .A2(n23262), .ZN(n23812) );
  OR3_X1 U18461 ( .A1(n25398), .A2(n26070), .A3(net714551), .ZN(n23810) );
  AOI21_X1 U18462 ( .B1(n23979), .B2(n24348), .A(n24538), .ZN(n23809) );
  NOR2_X1 U18463 ( .A1(n23813), .A2(net715598), .ZN(n26100) );
  OAI22_X1 U18464 ( .A1(n1692), .A2(net718432), .B1(net715420), .B2(net741572), 
        .ZN(n23813) );
  OR2_X1 U18465 ( .A1(n23814), .A2(n26068), .ZN(net766153) );
  AOI21_X1 U18466 ( .B1(net746753), .B2(n24351), .A(n23815), .ZN(n23814) );
  NAND3_X1 U18467 ( .A1(net714845), .A2(n24361), .A3(n23973), .ZN(n23815) );
  NAND3_X1 U18468 ( .A1(n23816), .A2(n23817), .A3(n23818), .ZN(n26106) );
  NAND2_X1 U18469 ( .A1(n25390), .A2(n14758), .ZN(n23818) );
  NAND2_X1 U18470 ( .A1(net718341), .A2(n24784), .ZN(n23817) );
  AOI22_X1 U18471 ( .A1(net715443), .A2(\core_inst/MEMWB_ALUOUT/DFF_28/N3 ), 
        .B1(net762717), .B2(n522), .ZN(n23816) );
  CLKBUF_X1 U18472 ( .A(net715445), .Z(net762717) );
  NAND2_X1 U18473 ( .A1(n23819), .A2(n26185), .ZN(n25511) );
  XNOR2_X1 U18474 ( .A(n23820), .B(net716215), .ZN(n23819) );
  NOR2_X1 U18475 ( .A1(n24323), .A2(n24125), .ZN(n23820) );
  OAI22_X1 U18476 ( .A1(n4352), .A2(net737101), .B1(net718133), .B2(net741306), 
        .ZN(net737937) );
  OR2_X2 U18477 ( .A1(n23821), .A2(n24125), .ZN(n24271) );
  NAND3_X1 U18478 ( .A1(n25508), .A2(n23822), .A3(n25416), .ZN(n23821) );
  OR2_X1 U18479 ( .A1(n25509), .A2(n23993), .ZN(n23822) );
  OAI21_X1 U18480 ( .B1(n24354), .B2(n26118), .A(n23823), .ZN(net714599) );
  NOR2_X1 U18481 ( .A1(n24541), .A2(n24200), .ZN(n23823) );
  NAND2_X1 U18482 ( .A1(n25942), .A2(n25981), .ZN(net714709) );
  AND2_X2 U18483 ( .A1(n23824), .A2(net755733), .ZN(net730300) );
  NOR2_X1 U18484 ( .A1(n24541), .A2(n24032), .ZN(n23824) );
  AND2_X2 U18485 ( .A1(n23825), .A2(n26021), .ZN(net755733) );
  NAND2_X1 U18486 ( .A1(net713627), .A2(n23826), .ZN(n23825) );
  XNOR2_X1 U18487 ( .A(n26201), .B(net716221), .ZN(n23826) );
  NOR3_X1 U18488 ( .A1(n23827), .A2(n23828), .A3(n23829), .ZN(net742224) );
  NOR2_X1 U18489 ( .A1(net742223), .A2(n25310), .ZN(n23829) );
  NOR2_X1 U18490 ( .A1(net718432), .A2(n1714), .ZN(n23828) );
  OAI22_X1 U18491 ( .A1(net786841), .A2(n4325), .B1(net742209), .B2(n25360), 
        .ZN(n23827) );
  OAI22_X1 U18492 ( .A1(net715421), .A2(n25362), .B1(net717718), .B2(n4346), 
        .ZN(net715575) );
  AOI21_X1 U18493 ( .B1(n23830), .B2(net758644), .A(net767320), .ZN(n25398) );
  NOR2_X1 U18494 ( .A1(n23831), .A2(net714855), .ZN(n23830) );
  NOR2_X1 U18495 ( .A1(n25824), .A2(n25825), .ZN(n23831) );
  OAI21_X1 U18496 ( .B1(n24176), .B2(n26034), .A(n23833), .ZN(net733283) );
  NOR2_X1 U18497 ( .A1(n23832), .A2(n24324), .ZN(n23833) );
  NAND2_X1 U18498 ( .A1(n23834), .A2(n23835), .ZN(net733282) );
  AND2_X1 U18499 ( .A1(n23832), .A2(n23837), .ZN(n23835) );
  INV_X1 U18500 ( .A(n24176), .ZN(n23837) );
  NAND2_X1 U18501 ( .A1(n26034), .A2(n23836), .ZN(n23834) );
  INV_X1 U18502 ( .A(n24324), .ZN(n23836) );
  NOR2_X1 U18503 ( .A1(n23838), .A2(n23850), .ZN(n26529) );
  OR2_X1 U18504 ( .A1(n23839), .A2(n23840), .ZN(n23850) );
  OAI21_X1 U18505 ( .B1(n23841), .B2(n23851), .A(net717091), .ZN(n23840) );
  AOI21_X1 U18506 ( .B1(n23842), .B2(n25935), .A(n23843), .ZN(n23839) );
  MUX2_X1 U18507 ( .A(n23844), .B(n23845), .S(n23846), .Z(n23838) );
  NOR3_X1 U18508 ( .A1(net714770), .A2(n25934), .A3(n23847), .ZN(n23846) );
  INV_X1 U18509 ( .A(n25397), .ZN(n23847) );
  INV_X1 U18510 ( .A(n23843), .ZN(n23845) );
  NAND2_X1 U18511 ( .A1(n23841), .A2(n23851), .ZN(n23843) );
  BUF_X1 U18512 ( .A(n25936), .Z(n23851) );
  NOR3_X1 U18513 ( .A1(n23848), .A2(n23849), .A3(n23841), .ZN(n23844) );
  NAND2_X1 U18514 ( .A1(n25940), .A2(n24288), .ZN(n23841) );
  INV_X1 U18515 ( .A(n25935), .ZN(n23849) );
  INV_X1 U18516 ( .A(n23842), .ZN(n23848) );
  NAND2_X1 U18517 ( .A1(n25437), .A2(n24568), .ZN(n23842) );
  NOR2_X1 U18518 ( .A1(n23853), .A2(n23852), .ZN(net715176) );
  OAI22_X1 U18519 ( .A1(net717106), .A2(n1714), .B1(net714943), .B2(n25310), 
        .ZN(n23852) );
  NOR2_X1 U18520 ( .A1(n4325), .A2(net750086), .ZN(n23853) );
  AOI21_X1 U18521 ( .B1(n23855), .B2(n23856), .A(n24196), .ZN(net729284) );
  NOR2_X1 U18522 ( .A1(net714096), .A2(n23857), .ZN(n23856) );
  NOR2_X1 U18523 ( .A1(n24191), .A2(n23854), .ZN(n23857) );
  NAND2_X1 U18524 ( .A1(n23858), .A2(n23859), .ZN(n23855) );
  INV_X1 U18525 ( .A(n23854), .ZN(n23859) );
  NAND2_X1 U18526 ( .A1(net714104), .A2(n26074), .ZN(n23858) );
  NOR2_X1 U18527 ( .A1(n23854), .A2(net717091), .ZN(net714096) );
  MUX2_X1 U18528 ( .A(net713892), .B(n26136), .S(n26076), .Z(n23854) );
  INV_X1 U18529 ( .A(net714749), .ZN(net714746) );
  NAND2_X1 U18530 ( .A1(n24268), .A2(n24608), .ZN(net713636) );
  NAND2_X1 U18531 ( .A1(n23861), .A2(n23860), .ZN(n25419) );
  AOI22_X1 U18532 ( .A1(net713679), .A2(net755207), .B1(net742324), .B2(n22673), .ZN(n23860) );
  AOI21_X1 U18533 ( .B1(net742315), .B2(n25788), .A(net755260), .ZN(n23861) );
  NAND2_X1 U18534 ( .A1(n23862), .A2(net89524), .ZN(net715795) );
  OAI211_X1 U18535 ( .C1(n11743), .C2(n25581), .A(net334510), .B(
        \core_inst/MEMWB_IR/DFF_30/N3 ), .ZN(n23862) );
  NOR2_X1 U18536 ( .A1(n23864), .A2(n23863), .ZN(net742068) );
  CLKBUF_X1 U18537 ( .A(n25369), .Z(n23863) );
  CLKBUF_X1 U18538 ( .A(n25368), .Z(n23864) );
  NOR2_X1 U18539 ( .A1(net715359), .A2(n23865), .ZN(n26062) );
  OR2_X1 U18540 ( .A1(net717543), .A2(net755207), .ZN(n23865) );
  NOR2_X1 U18541 ( .A1(n23866), .A2(n23867), .ZN(n24380) );
  XNOR2_X1 U18542 ( .A(n24336), .B(net718006), .ZN(n23867) );
  XNOR2_X1 U18543 ( .A(n24315), .B(n25589), .ZN(n23866) );
  OAI21_X1 U18544 ( .B1(n23868), .B2(n24566), .A(n23869), .ZN(n26173) );
  NOR2_X1 U18545 ( .A1(n23870), .A2(n23871), .ZN(n23869) );
  OAI22_X1 U18546 ( .A1(n24548), .A2(n24402), .B1(net750090), .B2(net755683), 
        .ZN(n23871) );
  OAI22_X1 U18547 ( .A1(net713707), .A2(net749902), .B1(net714871), .B2(
        net713683), .ZN(n23870) );
  NOR2_X1 U18548 ( .A1(n25792), .A2(n25791), .ZN(n23868) );
  NAND3_X1 U18549 ( .A1(n23873), .A2(n23872), .A3(n23874), .ZN(n26077) );
  NAND2_X1 U18550 ( .A1(n23875), .A2(net717876), .ZN(n23874) );
  AND2_X1 U18551 ( .A1(net737672), .A2(n25355), .ZN(n23875) );
  NAND2_X1 U18552 ( .A1(net718340), .A2(n24782), .ZN(n23873) );
  AOI22_X1 U18553 ( .A1(net715443), .A2(\core_inst/MEMWB_ALUOUT/DFF_13/N3 ), 
        .B1(net715445), .B2(n991), .ZN(n23872) );
  AND2_X1 U18554 ( .A1(n23978), .A2(net749410), .ZN(net755735) );
  NAND2_X1 U18555 ( .A1(n23876), .A2(net714756), .ZN(n25447) );
  NAND3_X1 U18556 ( .A1(net749930), .A2(n23877), .A3(n23878), .ZN(n23876) );
  OR2_X1 U18557 ( .A1(n25793), .A2(net713683), .ZN(n23878) );
  INV_X1 U18558 ( .A(n25795), .ZN(n23877) );
  NAND2_X1 U18559 ( .A1(n24380), .A2(n24381), .ZN(net715773) );
  NAND2_X1 U18560 ( .A1(net716385), .A2(n23879), .ZN(n26713) );
  AOI21_X1 U18561 ( .B1(n11848), .B2(n26573), .A(net712488), .ZN(n23879) );
  NAND2_X1 U18562 ( .A1(net714950), .A2(net714281), .ZN(n25939) );
  NOR2_X1 U18563 ( .A1(n23880), .A2(n23881), .ZN(n25776) );
  OAI22_X1 U18564 ( .A1(n25789), .A2(net734022), .B1(net762729), .B2(net714494), .ZN(n23881) );
  OAI22_X1 U18565 ( .A1(n26064), .A2(net780556), .B1(n24276), .B2(n26071), 
        .ZN(n23880) );
  NAND2_X1 U18566 ( .A1(net716385), .A2(n23882), .ZN(n26716) );
  AOI21_X1 U18567 ( .B1(n5577), .B2(n26459), .A(n26574), .ZN(n23882) );
  NOR2_X1 U18568 ( .A1(n23883), .A2(net713154), .ZN(n25383) );
  XNOR2_X1 U18569 ( .A(n23884), .B(n23885), .ZN(n23883) );
  XNOR2_X1 U18570 ( .A(n23892), .B(n24278), .ZN(n23885) );
  CLKBUF_X1 U18571 ( .A(n24029), .Z(n23892) );
  OAI21_X1 U18572 ( .B1(n26069), .B2(n23891), .A(n23886), .ZN(n23884) );
  AOI21_X1 U18573 ( .B1(n23887), .B2(n24549), .A(n23888), .ZN(n23886) );
  NAND2_X1 U18574 ( .A1(net714164), .A2(n23889), .ZN(n23887) );
  INV_X1 U18575 ( .A(n24317), .ZN(n23889) );
  OR2_X1 U18576 ( .A1(net714157), .A2(n23890), .ZN(n23891) );
  NAND2_X1 U18577 ( .A1(net742326), .A2(n24549), .ZN(n23890) );
  NAND2_X1 U18578 ( .A1(n23893), .A2(net749930), .ZN(n25379) );
  NOR2_X1 U18579 ( .A1(n25513), .A2(n25795), .ZN(n23893) );
  AND2_X1 U18580 ( .A1(net714754), .A2(n23894), .ZN(n26069) );
  NAND2_X1 U18581 ( .A1(n23895), .A2(n23896), .ZN(n23894) );
  NAND2_X1 U18582 ( .A1(n25379), .A2(net749558), .ZN(n23895) );
  CLKBUF_X1 U18583 ( .A(net714756), .Z(net749558) );
  AND2_X1 U18584 ( .A1(n26131), .A2(n23897), .ZN(net758890) );
  NOR2_X1 U18585 ( .A1(n24551), .A2(n25513), .ZN(n23897) );
  NAND2_X1 U18586 ( .A1(n23898), .A2(n25831), .ZN(n26181) );
  NOR2_X1 U18587 ( .A1(n25830), .A2(n25829), .ZN(n23898) );
  INV_X1 U18588 ( .A(n23899), .ZN(n25831) );
  OAI22_X1 U18589 ( .A1(net765629), .A2(n1187), .B1(net741958), .B2(n4415), 
        .ZN(n23899) );
  AOI21_X1 U18590 ( .B1(n24351), .B2(net746753), .A(n23900), .ZN(n24403) );
  NAND3_X1 U18591 ( .A1(net749798), .A2(n23973), .A3(net714845), .ZN(n23900)
         );
  NAND2_X1 U18592 ( .A1(n23909), .A2(net714529), .ZN(net714531) );
  INV_X1 U18593 ( .A(net714539), .ZN(net714547) );
  AOI21_X1 U18594 ( .B1(net742061), .B2(net714533), .A(n23901), .ZN(net714532)
         );
  NAND3_X1 U18595 ( .A1(n23902), .A2(n23903), .A3(n23904), .ZN(n23901) );
  NAND4_X1 U18596 ( .A1(n23905), .A2(net712872), .A3(n24319), .A4(net714539), 
        .ZN(n23904) );
  INV_X1 U18597 ( .A(n23906), .ZN(n23905) );
  NAND2_X1 U18598 ( .A1(n24335), .A2(net762673), .ZN(n23906) );
  AOI21_X1 U18599 ( .B1(n23907), .B2(net714539), .A(net713154), .ZN(n23903) );
  OAI21_X1 U18600 ( .B1(net714542), .B2(n23908), .A(net713923), .ZN(n23907) );
  NAND2_X1 U18601 ( .A1(n24089), .A2(net762673), .ZN(n23908) );
  INV_X1 U18602 ( .A(net713924), .ZN(net762673) );
  OAI21_X1 U18603 ( .B1(net712880), .B2(net713924), .A(net714545), .ZN(n23902)
         );
  INV_X1 U18604 ( .A(net714530), .ZN(net714533) );
  NAND2_X1 U18605 ( .A1(net718400), .A2(net714545), .ZN(net714530) );
  NAND2_X1 U18606 ( .A1(n24094), .A2(n25992), .ZN(net714539) );
  NAND2_X1 U18607 ( .A1(n25424), .A2(n23910), .ZN(net714529) );
  AND2_X1 U18608 ( .A1(n26404), .A2(net740526), .ZN(n23910) );
  NAND3_X1 U18609 ( .A1(n23911), .A2(net740493), .A3(n23912), .ZN(net740492)
         );
  INV_X1 U18610 ( .A(n25368), .ZN(n23912) );
  INV_X1 U18611 ( .A(n25369), .ZN(n23911) );
  NAND3_X1 U18612 ( .A1(n23913), .A2(net717843), .A3(n23915), .ZN(net715700)
         );
  AND3_X1 U18613 ( .A1(n25751), .A2(net715705), .A3(n23914), .ZN(n23915) );
  MUX2_X1 U18614 ( .A(net715706), .B(net715707), .S(s_MEMWB_IR[27]), .Z(n23914) );
  NOR2_X1 U18615 ( .A1(net740492), .A2(net749843), .ZN(n23913) );
  NAND4_X1 U18616 ( .A1(n23916), .A2(n23917), .A3(n23918), .A4(n23919), .ZN(
        n25368) );
  XNOR2_X1 U18617 ( .A(n1666), .B(n25584), .ZN(n23919) );
  XNOR2_X1 U18618 ( .A(n1665), .B(n25583), .ZN(n23918) );
  XNOR2_X1 U18619 ( .A(n25593), .B(net717830), .ZN(n23917) );
  XNOR2_X1 U18620 ( .A(net717952), .B(n25591), .ZN(n23916) );
  NAND2_X1 U18621 ( .A1(net713468), .A2(n26041), .ZN(n23920) );
  INV_X1 U18622 ( .A(n23921), .ZN(n24395) );
  OAI22_X1 U18623 ( .A1(net718134), .A2(n1655), .B1(n25595), .B2(n4412), .ZN(
        n23921) );
  MUX2_X1 U18624 ( .A(n23947), .B(n24262), .S(n25748), .Z(net762761) );
  INV_X1 U18625 ( .A(net740492), .ZN(net715669) );
  NOR2_X1 U18626 ( .A1(n23922), .A2(n23923), .ZN(n24136) );
  OAI22_X1 U18627 ( .A1(n1708), .A2(net715419), .B1(net742223), .B2(n25348), 
        .ZN(n23923) );
  OAI22_X1 U18628 ( .A1(net715421), .A2(n25361), .B1(net749443), .B2(n4397), 
        .ZN(n23922) );
  INV_X1 U18629 ( .A(n23924), .ZN(n26222) );
  MUX2_X1 U18630 ( .A(n24136), .B(n5585), .S(net741686), .Z(n23924) );
  NAND2_X1 U18631 ( .A1(n24544), .A2(n25788), .ZN(n23925) );
  AOI22_X1 U18632 ( .A1(n22673), .A2(net767330), .B1(net755207), .B2(net713681), .ZN(n23926) );
  NAND3_X1 U18633 ( .A1(n23926), .A2(n24558), .A3(n23925), .ZN(n24524) );
  AND2_X2 U18634 ( .A1(n23928), .A2(n23929), .ZN(n24033) );
  NAND2_X1 U18635 ( .A1(n23927), .A2(net787518), .ZN(n23929) );
  NOR2_X1 U18636 ( .A1(n25764), .A2(n25763), .ZN(n23927) );
  NAND2_X1 U18637 ( .A1(net741686), .A2(n17743), .ZN(n23928) );
  INV_X1 U18638 ( .A(net714948), .ZN(net714610) );
  AOI21_X1 U18639 ( .B1(n23930), .B2(n23948), .A(n25394), .ZN(net714948) );
  NOR2_X1 U18640 ( .A1(n24029), .A2(n24265), .ZN(n23930) );
  AOI21_X1 U18641 ( .B1(n23931), .B2(net714858), .A(n24040), .ZN(net714975) );
  NAND2_X1 U18642 ( .A1(n25828), .A2(n24575), .ZN(n23931) );
  NAND3_X1 U18643 ( .A1(n23932), .A2(n25385), .A3(n25386), .ZN(n24039) );
  AOI21_X1 U18644 ( .B1(net749274), .B2(net365821), .A(n25387), .ZN(n23932) );
  NOR2_X1 U18645 ( .A1(n25828), .A2(net767335), .ZN(n24040) );
  XNOR2_X1 U18646 ( .A(n24039), .B(net716223), .ZN(n23933) );
  MUX2_X1 U18647 ( .A(n23947), .B(n24262), .S(n25748), .Z(n23934) );
  AOI21_X1 U18648 ( .B1(net740075), .B2(net715666), .A(net718033), .ZN(
        net765400) );
  NOR2_X1 U18649 ( .A1(n23935), .A2(net767320), .ZN(net714754) );
  OAI21_X1 U18650 ( .B1(net742146), .B2(net755139), .A(net714860), .ZN(n23935)
         );
  NAND2_X1 U18651 ( .A1(n23937), .A2(n23936), .ZN(net738839) );
  NAND2_X1 U18652 ( .A1(net724913), .A2(n24351), .ZN(n23936) );
  INV_X1 U18653 ( .A(net714122), .ZN(net724913) );
  NOR2_X1 U18654 ( .A1(net714770), .A2(n25427), .ZN(n23937) );
  XNOR2_X1 U18655 ( .A(n24347), .B(net742324), .ZN(net724910) );
  INV_X1 U18656 ( .A(n23939), .ZN(n23938) );
  OAI21_X1 U18657 ( .B1(n26572), .B2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [8]), .A(n26576), .ZN(n23939) );
  NAND2_X1 U18658 ( .A1(net716385), .A2(n23940), .ZN(n26707) );
  AOI21_X1 U18659 ( .B1(n6460), .B2(n26576), .A(n26575), .ZN(n23940) );
  AOI21_X1 U18660 ( .B1(net749363), .B2(n23941), .A(n25749), .ZN(net773961) );
  NOR3_X1 U18661 ( .A1(net717843), .A2(n25748), .A3(n25750), .ZN(net773962) );
  OAI211_X1 U18662 ( .C1(n23942), .C2(n1684), .A(net713480), .B(n22742), .ZN(
        \core_inst/IDEX_RF_ADDR_DEST/DFF_4/N3 ) );
  NAND2_X1 U18663 ( .A1(net765341), .A2(n18136), .ZN(n23942) );
  OAI211_X1 U18664 ( .C1(n25747), .C2(n24316), .A(n24135), .B(
        \cu_inst/FW_UNIT/ITD_EXMEM/N14 ), .ZN(net750145) );
  AND2_X1 U18666 ( .A1(n24535), .A2(n24261), .ZN(n23944) );
  NAND2_X1 U18667 ( .A1(net717742), .A2(n24038), .ZN(net717760) );
  NAND2_X1 U18668 ( .A1(net717742), .A2(net715647), .ZN(n25595) );
  AND2_X1 U18669 ( .A1(net715672), .A2(net717742), .ZN(n24569) );
  AND2_X1 U18670 ( .A1(net717742), .A2(n24360), .ZN(net732533) );
  AND2_X1 U18671 ( .A1(net717742), .A2(n24038), .ZN(n24320) );
  CLKBUF_X1 U18672 ( .A(net717742), .Z(net749922) );
  BUF_X1 U18673 ( .A(net717760), .Z(net762680) );
  BUF_X1 U18674 ( .A(net717760), .Z(net750085) );
  BUF_X1 U18675 ( .A(net717760), .Z(net750086) );
  NAND2_X1 U18676 ( .A1(net715176), .A2(net715175), .ZN(net713710) );
  OR2_X1 U18677 ( .A1(n24088), .A2(n24033), .ZN(n23948) );
  OAI21_X1 U18678 ( .B1(n23949), .B2(net714610), .A(net730300), .ZN(n23950) );
  AOI211_X1 U18679 ( .C1(n24339), .C2(n24034), .A(n23949), .B(net750290), .ZN(
        n26020) );
  NAND3_X1 U18680 ( .A1(net728823), .A2(net728824), .A3(net769908), .ZN(n25397) );
  INV_X1 U18681 ( .A(net714756), .ZN(net769908) );
  AND3_X1 U18682 ( .A1(n23950), .A2(net749338), .A3(net749905), .ZN(n24139) );
  AOI21_X1 U18683 ( .B1(n24139), .B2(net738443), .A(net713167), .ZN(n23951) );
  INV_X1 U18684 ( .A(n23951), .ZN(n23957) );
  AOI21_X1 U18685 ( .B1(net765361), .B2(n23958), .A(n23959), .ZN(net713803) );
  INV_X1 U18686 ( .A(net765361), .ZN(net713813) );
  OAI22_X1 U18687 ( .A1(net742209), .A2(n25364), .B1(net717718), .B2(n4394), 
        .ZN(n25764) );
  XNOR2_X1 U18688 ( .A(n25585), .B(net366479), .ZN(n24281) );
  NOR2_X1 U18689 ( .A1(net713677), .A2(n24281), .ZN(n25825) );
  XNOR2_X1 U18690 ( .A(n26198), .B(net716215), .ZN(n23952) );
  AOI21_X1 U18691 ( .B1(n25824), .B2(net714977), .A(n25825), .ZN(net714756) );
  NAND2_X1 U18692 ( .A1(n25827), .A2(n25826), .ZN(n23972) );
  XNOR2_X1 U18693 ( .A(n23972), .B(net716221), .ZN(n24124) );
  NAND2_X1 U18694 ( .A1(n24124), .A2(net731329), .ZN(net715032) );
  NAND2_X1 U18695 ( .A1(n25837), .A2(n25836), .ZN(n25903) );
  XNOR2_X1 U18696 ( .A(n25903), .B(net716215), .ZN(n25845) );
  OR2_X2 U18697 ( .A1(n25845), .A2(n26212), .ZN(n25935) );
  NAND2_X1 U18698 ( .A1(n24350), .A2(n25935), .ZN(net714751) );
  AND3_X1 U18699 ( .A1(n26564), .A2(n24528), .A3(n25943), .ZN(net712879) );
  OAI21_X1 U18700 ( .B1(n23953), .B2(n26705), .A(n22874), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_18/N3 ) );
  MUX2_X1 U18701 ( .A(n26088), .B(n5587), .S(net741686), .Z(n23970) );
  NAND2_X1 U18702 ( .A1(n25844), .A2(n25843), .ZN(n24280) );
  XNOR2_X1 U18703 ( .A(n24280), .B(net366479), .ZN(n24302) );
  NAND2_X1 U18704 ( .A1(n24302), .A2(n24547), .ZN(n24197) );
  NAND2_X1 U18705 ( .A1(n25846), .A2(n26067), .ZN(net714612) );
  MUX2_X1 U18706 ( .A(n17924), .B(n25392), .S(net787526), .Z(net767335) );
  OAI21_X1 U18707 ( .B1(n25366), .B2(n26130), .A(n22868), .ZN(n23964) );
  OAI21_X1 U18708 ( .B1(n23964), .B2(net749936), .A(net713829), .ZN(n23963) );
  NAND2_X1 U18709 ( .A1(n25422), .A2(n26139), .ZN(n23962) );
  NAND3_X1 U18710 ( .A1(n26141), .A2(n26139), .A3(n24142), .ZN(n23960) );
  INV_X1 U18711 ( .A(n26142), .ZN(n23965) );
  NAND4_X1 U18712 ( .A1(n26142), .A2(net713810), .A3(n24096), .A4(n24282), 
        .ZN(n23954) );
  NOR2_X1 U18713 ( .A1(n24297), .A2(n26138), .ZN(n23958) );
  NOR2_X1 U18714 ( .A1(n25422), .A2(n23965), .ZN(n23955) );
  NAND3_X1 U18715 ( .A1(n23957), .A2(n26141), .A3(n24142), .ZN(n23956) );
  NOR2_X1 U18716 ( .A1(n23954), .A2(net712880), .ZN(net713805) );
  OAI211_X1 U18717 ( .C1(net749400), .C2(n24297), .A(n23956), .B(n23955), .ZN(
        net713804) );
  BUF_X1 U18718 ( .A(n26042), .Z(n24547) );
  MUX2_X1 U18719 ( .A(n26112), .B(\core_inst/EXMEM_NPC/DFF_6/N3 ), .S(
        net741686), .Z(net767357) );
  BUF_X1 U18720 ( .A(n24137), .Z(n24572) );
  CLKBUF_X1 U18721 ( .A(net780598), .Z(net767352) );
  AND2_X1 U18722 ( .A1(n25837), .A2(n25836), .ZN(n23966) );
  CLKBUF_X1 U18723 ( .A(n25887), .Z(n23967) );
  INV_X1 U18724 ( .A(net762579), .ZN(net767341) );
  INV_X1 U18725 ( .A(net762579), .ZN(net718134) );
  CLKBUF_X1 U18726 ( .A(n25824), .Z(n23968) );
  AND2_X1 U18727 ( .A1(n25793), .A2(net749725), .ZN(n25824) );
  INV_X1 U18728 ( .A(net749832), .ZN(net767330) );
  MUX2_X1 U18729 ( .A(n26088), .B(n5587), .S(net741686), .Z(n23969) );
  CLKBUF_X1 U18730 ( .A(n26150), .Z(n24175) );
  OR2_X1 U18731 ( .A1(n24347), .A2(net742325), .ZN(n24351) );
  NAND2_X1 U18732 ( .A1(n25587), .A2(n24576), .ZN(n23973) );
  AND2_X1 U18733 ( .A1(n25848), .A2(n25847), .ZN(n23974) );
  CLKBUF_X1 U18734 ( .A(n24271), .Z(n23975) );
  NOR2_X1 U18735 ( .A1(net715221), .A2(n25821), .ZN(n23976) );
  XNOR2_X1 U18736 ( .A(net742241), .B(net716215), .ZN(n23977) );
  OR2_X1 U18737 ( .A1(net715528), .A2(net715586), .ZN(net718152) );
  AOI21_X1 U18738 ( .B1(n25898), .B2(n23977), .A(n24202), .ZN(n23978) );
  INV_X2 U18739 ( .A(net755610), .ZN(net748269) );
  MUX2_X1 U18740 ( .A(\core_inst/EXMEM_NPC/DFF_4/N3 ), .B(n26096), .S(
        net787528), .Z(n24192) );
  BUF_X2 U18741 ( .A(n26022), .Z(n24300) );
  CLKBUF_X3 U18742 ( .A(net749312), .Z(net718367) );
  INV_X2 U18743 ( .A(net718367), .ZN(net739078) );
  BUF_X2 U18744 ( .A(n26134), .Z(n24233) );
  BUF_X2 U18745 ( .A(n26134), .Z(n24270) );
  BUF_X2 U18746 ( .A(net717060), .Z(net762753) );
  NOR2_X1 U18747 ( .A1(net714602), .A2(n25834), .ZN(n26564) );
  AND2_X1 U18748 ( .A1(net765341), .A2(n26559), .ZN(n23980) );
  AND2_X1 U18749 ( .A1(net742576), .A2(n26458), .ZN(n23982) );
  AND2_X1 U18750 ( .A1(net742576), .A2(net712808), .ZN(n23983) );
  AND2_X1 U18751 ( .A1(net716243), .A2(n26534), .ZN(n23985) );
  AND2_X1 U18752 ( .A1(net742648), .A2(n26530), .ZN(n23986) );
  AND2_X1 U18753 ( .A1(net742649), .A2(net713438), .ZN(n23987) );
  AND2_X1 U18754 ( .A1(net785255), .A2(n26568), .ZN(n23988) );
  AND2_X1 U18755 ( .A1(net742648), .A2(n26410), .ZN(n23989) );
  AND2_X1 U18756 ( .A1(net760161), .A2(n24168), .ZN(n23990) );
  BUF_X1 U18757 ( .A(n24329), .Z(n26031) );
  BUF_X1 U18758 ( .A(net713906), .Z(net742259) );
  INV_X1 U18759 ( .A(net755139), .ZN(net749612) );
  INV_X1 U18760 ( .A(n25989), .ZN(n24158) );
  INV_X2 U18761 ( .A(n24004), .ZN(n20351) );
  INV_X2 U18762 ( .A(n24005), .ZN(n20368) );
  INV_X2 U18763 ( .A(n24006), .ZN(n20334) );
  INV_X2 U18764 ( .A(n24002), .ZN(n20394) );
  INV_X2 U18765 ( .A(n24003), .ZN(n20375) );
  INV_X2 U18766 ( .A(n24000), .ZN(n20521) );
  INV_X2 U18767 ( .A(n23997), .ZN(n20686) );
  INV_X2 U18768 ( .A(n23999), .ZN(n20549) );
  INV_X2 U18769 ( .A(n23998), .ZN(n20582) );
  INV_X2 U18770 ( .A(n23996), .ZN(n20502) );
  INV_X2 U18771 ( .A(n24001), .ZN(n20445) );
  BUF_X2 U18772 ( .A(n20547), .Z(n23999) );
  BUF_X2 U18773 ( .A(n20581), .Z(n23998) );
  BUF_X2 U18774 ( .A(n20519), .Z(n24000) );
  BUF_X2 U18775 ( .A(n20684), .Z(n23997) );
  BUF_X2 U18776 ( .A(n20367), .Z(n24005) );
  BUF_X2 U18777 ( .A(n20373), .Z(n24003) );
  BUF_X2 U18778 ( .A(n20392), .Z(n24002) );
  BUF_X2 U18779 ( .A(n20443), .Z(n24001) );
  BUF_X2 U18780 ( .A(n20501), .Z(n23996) );
  BUF_X2 U18781 ( .A(n20350), .Z(n24004) );
  BUF_X2 U18782 ( .A(n20333), .Z(n24006) );
  NOR2_X1 U18783 ( .A1(n20154), .A2(n20220), .ZN(n20611) );
  NOR2_X1 U18784 ( .A1(n20200), .A2(n20372), .ZN(n20481) );
  NOR2_X1 U18785 ( .A1(n20260), .A2(n20431), .ZN(n20462) );
  NOR2_X1 U18786 ( .A1(n20200), .A2(n20332), .ZN(n20313) );
  NOR2_X1 U18787 ( .A1(n20220), .A2(n20293), .ZN(n20294) );
  NOR2_X1 U18788 ( .A1(n20200), .A2(n20260), .ZN(n20241) );
  NOR2_X1 U18789 ( .A1(n20200), .A2(n20240), .ZN(n20221) );
  NOR2_X1 U18790 ( .A1(n20200), .A2(n20220), .ZN(n20202) );
  NOR2_X1 U18791 ( .A1(n20154), .A2(n20332), .ZN(n20667) );
  NOR2_X1 U18792 ( .A1(n20154), .A2(n20260), .ZN(n20650) );
  NOR2_X1 U18793 ( .A1(n20154), .A2(n20240), .ZN(n20630) );
  NOR2_X1 U18794 ( .A1(n20154), .A2(n20201), .ZN(n20592) );
  NOR2_X1 U18795 ( .A1(n20220), .A2(n20431), .ZN(n20432) );
  NOR2_X1 U18796 ( .A1(n20201), .A2(n20431), .ZN(n20398) );
  NOR2_X1 U18797 ( .A1(n20372), .A2(n20293), .ZN(n20370) );
  NOR2_X1 U18798 ( .A1(n20201), .A2(n20293), .ZN(n20261) );
  NOR2_X1 U18799 ( .A1(n20153), .A2(n20200), .ZN(n20704) );
  INV_X2 U18800 ( .A(n24614), .ZN(n23994) );
  BUF_X1 U18801 ( .A(n19334), .Z(n24007) );
  BUF_X1 U18802 ( .A(n18329), .Z(net767214) );
  INV_X2 U18803 ( .A(n24613), .ZN(n23995) );
  INV_X1 U18804 ( .A(net713728), .ZN(net767234) );
  INV_X1 U18805 ( .A(n26606), .ZN(n26608) );
  AND2_X1 U18806 ( .A1(net714657), .A2(net714306), .ZN(n25893) );
  AND2_X1 U18807 ( .A1(net713966), .A2(net714934), .ZN(net735179) );
  INV_X1 U18808 ( .A(n25860), .ZN(n24245) );
  INV_X1 U18809 ( .A(net749894), .ZN(net713767) );
  BUF_X1 U18810 ( .A(n26027), .Z(n24536) );
  AND2_X1 U18811 ( .A1(net737713), .A2(net713863), .ZN(net749894) );
  AND2_X1 U18812 ( .A1(n25579), .A2(net713863), .ZN(n26056) );
  INV_X1 U18813 ( .A(n26182), .ZN(n24371) );
  INV_X1 U18814 ( .A(net714275), .ZN(net714182) );
  INV_X1 U18815 ( .A(net713985), .ZN(net742087) );
  MUX2_X1 U18816 ( .A(n17743), .B(n24092), .S(net716237), .Z(n24341) );
  INV_X1 U18817 ( .A(n26080), .ZN(n26081) );
  INV_X1 U18818 ( .A(n26717), .ZN(n24008) );
  AND2_X1 U18819 ( .A1(net713412), .A2(net713414), .ZN(n26717) );
  INV_X2 U18820 ( .A(n20221), .ZN(n20223) );
  INV_X2 U18821 ( .A(n20462), .ZN(n20464) );
  INV_X2 U18822 ( .A(n20202), .ZN(n20204) );
  INV_X2 U18823 ( .A(n20241), .ZN(n20243) );
  INV_X2 U18824 ( .A(n20667), .ZN(n20668) );
  INV_X2 U18825 ( .A(n20481), .ZN(n20483) );
  INV_X2 U18826 ( .A(n20704), .ZN(n20706) );
  INV_X2 U18827 ( .A(n20294), .ZN(n20296) );
  INV_X2 U18828 ( .A(n20313), .ZN(n20315) );
  INV_X2 U18829 ( .A(n20611), .ZN(n20613) );
  INV_X2 U18830 ( .A(n20630), .ZN(n20632) );
  INV_X2 U18831 ( .A(n20261), .ZN(n20263) );
  INV_X2 U18832 ( .A(n20432), .ZN(n20433) );
  INV_X2 U18833 ( .A(n20370), .ZN(n20371) );
  INV_X2 U18834 ( .A(n20592), .ZN(n20593) );
  INV_X2 U18835 ( .A(n20398), .ZN(n20400) );
  INV_X2 U18836 ( .A(n20650), .ZN(n20651) );
  BUF_X2 U18837 ( .A(n20261), .Z(n24025) );
  AOI211_X1 U18838 ( .C1(net767173), .C2(n534), .A(n24482), .B(n24483), .ZN(
        n24470) );
  BUF_X2 U18839 ( .A(n20704), .Z(n24023) );
  BUF_X2 U18840 ( .A(n20630), .Z(n24024) );
  BUF_X2 U18841 ( .A(n20611), .Z(n24022) );
  BUF_X2 U18842 ( .A(n20481), .Z(n24021) );
  BUF_X2 U18843 ( .A(n20462), .Z(n24020) );
  BUF_X2 U18844 ( .A(n20313), .Z(n24019) );
  BUF_X2 U18845 ( .A(n20294), .Z(n24018) );
  BUF_X2 U18846 ( .A(n20241), .Z(n24017) );
  BUF_X2 U18847 ( .A(n20221), .Z(n24016) );
  BUF_X2 U18848 ( .A(n20202), .Z(n24015) );
  BUF_X2 U18849 ( .A(n20667), .Z(n24014) );
  BUF_X2 U18850 ( .A(n20650), .Z(n24013) );
  BUF_X2 U18851 ( .A(n20592), .Z(n24012) );
  NAND2_X1 U18852 ( .A1(net767171), .A2(n23261), .ZN(n24505) );
  AOI21_X1 U18853 ( .B1(net767167), .B2(n956), .A(n24506), .ZN(n24504) );
  AOI211_X1 U18854 ( .C1(net767173), .C2(n964), .A(n24517), .B(n24518), .ZN(
        n24513) );
  NAND2_X1 U18855 ( .A1(net767173), .A2(n23260), .ZN(n24052) );
  NOR2_X1 U18856 ( .A1(net767172), .A2(n2090), .ZN(n24064) );
  BUF_X2 U18857 ( .A(n20398), .Z(n24010) );
  BUF_X2 U18858 ( .A(n20370), .Z(n24009) );
  BUF_X2 U18859 ( .A(n20432), .Z(n24011) );
  INV_X2 U18860 ( .A(n26714), .ZN(n26715) );
  INV_X1 U18861 ( .A(n18347), .ZN(net767172) );
  INV_X1 U18862 ( .A(n18332), .ZN(net767171) );
  INV_X1 U18863 ( .A(n18398), .ZN(net767169) );
  INV_X1 U18864 ( .A(net713751), .ZN(net767221) );
  NOR2_X1 U18865 ( .A1(n26778), .A2(n20067), .ZN(n25667) );
  INV_X1 U18866 ( .A(n19294), .ZN(n26780) );
  NOR2_X2 U18867 ( .A1(s_WB_MUX_CONTROL[1]), .A2(s_WB_MUX_CONTROL[0]), .ZN(
        net712606) );
  INV_X1 U18868 ( .A(n26580), .ZN(n26581) );
  INV_X1 U18869 ( .A(n25580), .ZN(n26725) );
  AND2_X1 U18870 ( .A1(n26126), .A2(net713863), .ZN(net732750) );
  INV_X1 U18871 ( .A(n26011), .ZN(n26014) );
  INV_X1 U18872 ( .A(net714261), .ZN(net714240) );
  INV_X1 U18873 ( .A(n26154), .ZN(n26161) );
  INV_X1 U18874 ( .A(n26050), .ZN(n25996) );
  INV_X1 U18875 ( .A(n24379), .ZN(n26123) );
  INV_X1 U18876 ( .A(net713977), .ZN(net713869) );
  NOR2_X1 U18877 ( .A1(net712838), .A2(n6402), .ZN(n26457) );
  BUF_X1 U18878 ( .A(net728314), .Z(net755757) );
  INV_X1 U18879 ( .A(n26138), .ZN(n26139) );
  INV_X1 U18880 ( .A(n26010), .ZN(n26012) );
  OR2_X1 U18881 ( .A1(n24145), .A2(n24146), .ZN(net740679) );
  OAI21_X1 U18882 ( .B1(net749894), .B2(n24421), .A(n24422), .ZN(n24418) );
  INV_X1 U18883 ( .A(net714382), .ZN(net713874) );
  INV_X1 U18884 ( .A(n26053), .ZN(n26203) );
  AND2_X1 U18885 ( .A1(net732754), .A2(net767221), .ZN(net732762) );
  AND2_X1 U18886 ( .A1(n24088), .A2(n24033), .ZN(n25394) );
  INV_X1 U18887 ( .A(net713950), .ZN(net713829) );
  INV_X1 U18888 ( .A(net749977), .ZN(net767211) );
  INV_X1 U18889 ( .A(net714306), .ZN(net767209) );
  INV_X1 U18890 ( .A(net714267), .ZN(net767208) );
  INV_X1 U18891 ( .A(n26183), .ZN(n24373) );
  INV_X1 U18892 ( .A(n26001), .ZN(n26228) );
  INV_X1 U18893 ( .A(n26234), .ZN(n26240) );
  MUX2_X1 U18894 ( .A(\core_inst/EXMEM_NPC/DFF_14/N3 ), .B(n26091), .S(
        net716237), .Z(n26212) );
  INV_X1 U18895 ( .A(net713985), .ZN(net767206) );
  AND2_X1 U18896 ( .A1(net712499), .A2(n26478), .ZN(n26479) );
  BUF_X1 U18897 ( .A(net717104), .Z(net717105) );
  AND2_X1 U18898 ( .A1(net717048), .A2(n26467), .ZN(n26468) );
  AND2_X1 U18899 ( .A1(n25665), .A2(n26684), .ZN(n26506) );
  BUF_X2 U18900 ( .A(net717104), .Z(net765744) );
  AND2_X1 U18901 ( .A1(net717048), .A2(n26400), .ZN(n26401) );
  INV_X1 U18902 ( .A(n26704), .ZN(n26637) );
  AND2_X1 U18903 ( .A1(net712499), .A2(n26658), .ZN(n26418) );
  AND2_X1 U18904 ( .A1(net712499), .A2(n26661), .ZN(n26590) );
  AND2_X1 U18905 ( .A1(n25665), .A2(n26670), .ZN(n26390) );
  AND2_X1 U18906 ( .A1(net717048), .A2(n26526), .ZN(n26310) );
  AND2_X1 U18907 ( .A1(net712397), .A2(n26490), .ZN(n26491) );
  AND2_X1 U18908 ( .A1(net717049), .A2(n26448), .ZN(n26321) );
  AND2_X1 U18909 ( .A1(net717049), .A2(n26648), .ZN(n26649) );
  AND2_X1 U18910 ( .A1(net712397), .A2(n26299), .ZN(n26300) );
  AND2_X1 U18911 ( .A1(net717049), .A2(n26714), .ZN(n26694) );
  AND3_X1 U18912 ( .A1(n26274), .A2(n20041), .A3(n26273), .ZN(net717048) );
  NOR4_X1 U18913 ( .A1(n24447), .A2(n24448), .A3(n24449), .A4(n24450), .ZN(
        n24446) );
  AND3_X1 U18914 ( .A1(n26274), .A2(n20041), .A3(n26273), .ZN(n25665) );
  INV_X1 U18915 ( .A(net717049), .ZN(net765730) );
  AND3_X1 U18916 ( .A1(n26274), .A2(n20041), .A3(n26273), .ZN(net712499) );
  INV_X1 U18917 ( .A(net742017), .ZN(net767205) );
  AOI22_X1 U18918 ( .A1(net717050), .A2(n26639), .B1(n26717), .B2(n24042), 
        .ZN(n24041) );
  NAND4_X1 U18919 ( .A1(n24043), .A2(n24044), .A3(n24045), .A4(n24046), .ZN(
        n24042) );
  AND4_X1 U18920 ( .A1(n24491), .A2(n24492), .A3(n24493), .A4(n24494), .ZN(
        n24490) );
  NAND4_X1 U18921 ( .A1(n24451), .A2(n24452), .A3(n24453), .A4(n24454), .ZN(
        n24450) );
  AND2_X1 U18922 ( .A1(net713412), .A2(net713414), .ZN(n25664) );
  INV_X1 U18923 ( .A(n24496), .ZN(n24492) );
  NOR2_X1 U18924 ( .A1(n24049), .A2(n24050), .ZN(n24044) );
  AND2_X1 U18925 ( .A1(n18929), .A2(n18928), .ZN(n24432) );
  AND2_X1 U18926 ( .A1(n18763), .A2(n18762), .ZN(n26653) );
  NOR2_X1 U18927 ( .A1(n24511), .A2(n24512), .ZN(n24488) );
  AND2_X1 U18928 ( .A1(n18736), .A2(n18735), .ZN(n24441) );
  NAND4_X1 U18929 ( .A1(n24470), .A2(n24471), .A3(n24472), .A4(n24473), .ZN(
        n24447) );
  OAI211_X1 U18930 ( .C1(n18332), .C2(n546), .A(n24464), .B(n24465), .ZN(
        n24448) );
  AND2_X1 U18931 ( .A1(n18709), .A2(n18708), .ZN(n25543) );
  INV_X1 U18932 ( .A(n24456), .ZN(n24452) );
  AND2_X1 U18933 ( .A1(n18570), .A2(n18569), .ZN(n26520) );
  AND4_X1 U18934 ( .A1(n19958), .A2(n19959), .A3(n19960), .A4(n19961), .ZN(
        n26664) );
  AND2_X1 U18935 ( .A1(n18790), .A2(n18789), .ZN(n26275) );
  AND2_X1 U18936 ( .A1(n18983), .A2(n18982), .ZN(n26345) );
  AND2_X1 U18937 ( .A1(n18628), .A2(n18627), .ZN(n25556) );
  AND2_X1 U18938 ( .A1(n18682), .A2(n18681), .ZN(n26430) );
  AND2_X1 U18939 ( .A1(n18844), .A2(n18843), .ZN(n25564) );
  AND2_X1 U18940 ( .A1(n19854), .A2(n19853), .ZN(n26393) );
  AND2_X1 U18941 ( .A1(n19722), .A2(n19721), .ZN(n26449) );
  AND2_X1 U18942 ( .A1(n19832), .A2(n19831), .ZN(n26632) );
  AND2_X1 U18943 ( .A1(n19700), .A2(n19699), .ZN(n26471) );
  AND2_X1 U18944 ( .A1(n19656), .A2(n19655), .ZN(n26460) );
  OAI211_X1 U18945 ( .C1(net767232), .C2(n979), .A(n24497), .B(n24498), .ZN(
        n24496) );
  NOR2_X1 U18946 ( .A1(n24500), .A2(n24501), .ZN(n24489) );
  NOR2_X1 U18947 ( .A1(n24047), .A2(n24048), .ZN(n24045) );
  OAI211_X1 U18948 ( .C1(n18401), .C2(n2081), .A(n24051), .B(n24052), .ZN(
        n24050) );
  NOR2_X1 U18949 ( .A1(n24063), .A2(n24064), .ZN(n24043) );
  AND2_X1 U18950 ( .A1(n19568), .A2(n19567), .ZN(n26583) );
  AND2_X1 U18951 ( .A1(n19523), .A2(n19522), .ZN(n26303) );
  AND2_X1 U18952 ( .A1(n19678), .A2(n19677), .ZN(n26411) );
  AND2_X1 U18953 ( .A1(n19612), .A2(n19611), .ZN(n26352) );
  NOR2_X1 U18954 ( .A1(n24475), .A2(n24476), .ZN(n24471) );
  AND2_X1 U18955 ( .A1(n19590), .A2(n19589), .ZN(n26383) );
  OAI211_X1 U18956 ( .C1(net767232), .C2(n549), .A(n24457), .B(n24458), .ZN(
        n24456) );
  AND2_X1 U18957 ( .A1(n19634), .A2(n19633), .ZN(n26329) );
  AND2_X1 U18958 ( .A1(n19876), .A2(n19875), .ZN(n26324) );
  AND2_X1 U18959 ( .A1(n19810), .A2(n19809), .ZN(n26421) );
  AND2_X1 U18960 ( .A1(n19037), .A2(n19036), .ZN(n26640) );
  INV_X1 U18961 ( .A(n25640), .ZN(n26670) );
  INV_X1 U18962 ( .A(n25630), .ZN(n26478) );
  AND3_X1 U18963 ( .A1(n18801), .A2(n18800), .A3(n18799), .ZN(n24837) );
  OAI22_X1 U18964 ( .A1(net767232), .A2(n24658), .B1(n2088), .B2(net716477), 
        .ZN(n24047) );
  AND3_X1 U18965 ( .A1(n18693), .A2(n18692), .A3(n18691), .ZN(n24839) );
  AND2_X1 U18966 ( .A1(n19919), .A2(n19918), .ZN(n25548) );
  AOI21_X1 U18967 ( .B1(net716461), .B2(n529), .A(n24455), .ZN(n24453) );
  AND3_X1 U18968 ( .A1(n18943), .A2(n24430), .A3(n24431), .ZN(n24433) );
  AND3_X1 U18969 ( .A1(n18639), .A2(n18638), .A3(n18637), .ZN(n24835) );
  AND3_X1 U18970 ( .A1(n18940), .A2(n18939), .A3(n18938), .ZN(n24434) );
  AND3_X1 U18971 ( .A1(n18747), .A2(n18746), .A3(n18745), .ZN(n24443) );
  AND3_X1 U18972 ( .A1(n20034), .A2(n20033), .A3(n20032), .ZN(n24075) );
  AND2_X1 U18973 ( .A1(n19120), .A2(n19119), .ZN(n26686) );
  AND3_X1 U18974 ( .A1(n18750), .A2(n24439), .A3(n24440), .ZN(n24442) );
  INV_X2 U18975 ( .A(n20155), .ZN(n25670) );
  INV_X1 U18976 ( .A(n25620), .ZN(n26706) );
  INV_X2 U18977 ( .A(n20183), .ZN(n25668) );
  NAND2_X1 U18978 ( .A1(n24480), .A2(n24481), .ZN(n24475) );
  AND2_X1 U18979 ( .A1(n19148), .A2(n19147), .ZN(n26291) );
  AND3_X1 U18980 ( .A1(n18804), .A2(n26277), .A3(n26276), .ZN(n25260) );
  AOI21_X1 U18981 ( .B1(n18312), .B2(n537), .A(n24474), .ZN(n24472) );
  AND3_X1 U18982 ( .A1(n19929), .A2(n19928), .A3(n19927), .ZN(n24834) );
  AND3_X1 U18983 ( .A1(n18777), .A2(n26655), .A3(n26654), .ZN(n25262) );
  AND3_X1 U18984 ( .A1(n18720), .A2(n18719), .A3(n18718), .ZN(n24833) );
  AND2_X1 U18985 ( .A1(n20024), .A2(n20023), .ZN(n24070) );
  INV_X1 U18986 ( .A(n25624), .ZN(n26669) );
  AND3_X1 U18987 ( .A1(n24466), .A2(n24467), .A3(n24468), .ZN(n24465) );
  INV_X1 U18988 ( .A(n24459), .ZN(n24457) );
  INV_X1 U18989 ( .A(n25638), .ZN(n26436) );
  AOI21_X1 U18990 ( .B1(n18312), .B2(n967), .A(n24516), .ZN(n24514) );
  AND3_X1 U18991 ( .A1(n18581), .A2(n18580), .A3(n18579), .ZN(n24840) );
  OAI22_X1 U18992 ( .A1(n18332), .A2(n24673), .B1(n24593), .B2(n18363), .ZN(
        n24063) );
  AND2_X1 U18993 ( .A1(n19898), .A2(n19897), .ZN(n24106) );
  AOI21_X1 U18994 ( .B1(n18307), .B2(n17790), .A(n24523), .ZN(n24519) );
  AND2_X1 U18995 ( .A1(n19235), .A2(n19234), .ZN(n26313) );
  NOR2_X1 U18996 ( .A1(n26272), .A2(n26271), .ZN(n26273) );
  AND2_X1 U18997 ( .A1(n20057), .A2(n20056), .ZN(n26439) );
  AND3_X1 U18998 ( .A1(n18855), .A2(n18854), .A3(n18853), .ZN(n24836) );
  AND2_X1 U18999 ( .A1(n19176), .A2(n19175), .ZN(n26374) );
  AND3_X1 U19000 ( .A1(n18994), .A2(n18993), .A3(n18992), .ZN(n24838) );
  AND2_X1 U19001 ( .A1(n19204), .A2(n19203), .ZN(n26482) );
  AOI21_X1 U19002 ( .B1(net716461), .B2(n959), .A(n24495), .ZN(n24493) );
  INV_X2 U19003 ( .A(n20134), .ZN(n25672) );
  INV_X1 U19004 ( .A(n25642), .ZN(n26661) );
  INV_X1 U19005 ( .A(n24499), .ZN(n24497) );
  AOI21_X1 U19006 ( .B1(n18306), .B2(n968), .A(n24522), .ZN(n24521) );
  AND3_X1 U19007 ( .A1(n18774), .A2(n18773), .A3(n18772), .ZN(n24841) );
  INV_X1 U19008 ( .A(n24053), .ZN(n24051) );
  AND2_X1 U19009 ( .A1(n19982), .A2(n19981), .ZN(n24080) );
  AND3_X1 U19010 ( .A1(n19908), .A2(n19907), .A3(n19906), .ZN(n24111) );
  INV_X1 U19011 ( .A(n25604), .ZN(n26490) );
  AND3_X1 U19012 ( .A1(n18997), .A2(n26347), .A3(n26346), .ZN(n25261) );
  OR4_X1 U19013 ( .A1(n25522), .A2(n25523), .A3(n19489), .A4(n19490), .ZN(
        n25518) );
  INV_X1 U19014 ( .A(n25606), .ZN(n26631) );
  AND3_X1 U19015 ( .A1(n19992), .A2(n19991), .A3(n19990), .ZN(n24085) );
  INV_X1 U19016 ( .A(n25648), .ZN(n26662) );
  NAND4_X1 U19017 ( .A1(n24502), .A2(n24503), .A3(n24504), .A4(n24505), .ZN(
        n24501) );
  INV_X1 U19018 ( .A(n25602), .ZN(n26448) );
  AND2_X1 U19019 ( .A1(n25722), .A2(n25721), .ZN(n26756) );
  INV_X1 U19020 ( .A(n25627), .ZN(n26652) );
  INV_X1 U19021 ( .A(n25656), .ZN(n26675) );
  INV_X1 U19022 ( .A(n25618), .ZN(n26400) );
  INV_X1 U19023 ( .A(n25616), .ZN(n26327) );
  INV_X1 U19024 ( .A(n25610), .ZN(n26600) );
  AND2_X1 U19025 ( .A1(n25691), .A2(n25690), .ZN(n26773) );
  AND2_X1 U19026 ( .A1(n25724), .A2(n25723), .ZN(n25641) );
  AND2_X1 U19027 ( .A1(n25691), .A2(n25690), .ZN(n25606) );
  AND2_X1 U19028 ( .A1(n25714), .A2(n25713), .ZN(n25631) );
  AND2_X1 U19029 ( .A1(n25691), .A2(n25690), .ZN(n25607) );
  AND2_X1 U19030 ( .A1(n25689), .A2(n25688), .ZN(n26774) );
  AND2_X1 U19031 ( .A1(n25724), .A2(n25723), .ZN(n26755) );
  BUF_X2 U19032 ( .A(n20155), .Z(n25671) );
  AND2_X1 U19033 ( .A1(n25714), .A2(n25713), .ZN(n26760) );
  AND2_X1 U19034 ( .A1(n25714), .A2(n25713), .ZN(n25630) );
  AND2_X1 U19035 ( .A1(n25689), .A2(n25688), .ZN(n25605) );
  AND2_X1 U19036 ( .A1(n25724), .A2(n25723), .ZN(n25640) );
  BUF_X2 U19037 ( .A(n20183), .Z(n25669) );
  AND2_X1 U19038 ( .A1(n25689), .A2(n25688), .ZN(n25604) );
  AND2_X1 U19039 ( .A1(n25722), .A2(n25721), .ZN(n25638) );
  AND2_X1 U19040 ( .A1(n25722), .A2(n25721), .ZN(n25639) );
  INV_X1 U19041 ( .A(n25634), .ZN(n26467) );
  AND2_X1 U19042 ( .A1(n25732), .A2(n25731), .ZN(n25648) );
  AND2_X1 U19043 ( .A1(n25732), .A2(n25731), .ZN(n26751) );
  INV_X1 U19044 ( .A(n25608), .ZN(n26299) );
  AND2_X1 U19045 ( .A1(net715892), .A2(n25708), .ZN(n25625) );
  INV_X1 U19046 ( .A(n26255), .ZN(n26510) );
  AND2_X1 U19047 ( .A1(net715892), .A2(n25708), .ZN(n25624) );
  AND2_X1 U19048 ( .A1(net715892), .A2(n25708), .ZN(n26764) );
  AND2_X1 U19049 ( .A1(n25726), .A2(n25725), .ZN(n26754) );
  INV_X1 U19050 ( .A(n25660), .ZN(n26684) );
  AND2_X1 U19051 ( .A1(n25726), .A2(n25725), .ZN(n25642) );
  INV_X1 U19052 ( .A(n25614), .ZN(n26648) );
  AND2_X1 U19053 ( .A1(n25726), .A2(n25725), .ZN(n25643) );
  BUF_X2 U19054 ( .A(n20134), .Z(n25673) );
  INV_X1 U19055 ( .A(n25650), .ZN(n26718) );
  INV_X1 U19056 ( .A(n25646), .ZN(n26526) );
  INV_X1 U19057 ( .A(n25644), .ZN(n26624) );
  INV_X1 U19058 ( .A(n25636), .ZN(n26603) );
  INV_X1 U19059 ( .A(n25654), .ZN(n26639) );
  INV_X1 U19060 ( .A(n26270), .ZN(n26272) );
  INV_X1 U19061 ( .A(n25652), .ZN(n26555) );
  AND2_X1 U19062 ( .A1(n25705), .A2(n25704), .ZN(n26766) );
  OAI22_X1 U19063 ( .A1(net767237), .A2(n24672), .B1(n2087), .B2(n18369), .ZN(
        n24053) );
  AND2_X1 U19064 ( .A1(n25705), .A2(n25704), .ZN(n25620) );
  INV_X1 U19065 ( .A(n25632), .ZN(n26658) );
  AND2_X1 U19066 ( .A1(n25705), .A2(n25704), .ZN(n25621) );
  AOI211_X1 U19067 ( .C1(net767239), .C2(n17926), .A(n24057), .B(n24058), .ZN(
        n24056) );
  AOI211_X1 U19068 ( .C1(n17936), .C2(net716405), .A(n24059), .B(n24060), .ZN(
        n24055) );
  AOI211_X1 U19069 ( .C1(net716417), .C2(n17927), .A(n24061), .B(n24062), .ZN(
        n24054) );
  INV_X1 U19070 ( .A(n24109), .ZN(n24108) );
  AND2_X1 U19071 ( .A1(n25687), .A2(n25686), .ZN(n26775) );
  AND2_X1 U19072 ( .A1(n25687), .A2(n25686), .ZN(n25602) );
  AND2_X1 U19073 ( .A1(n25687), .A2(n25686), .ZN(n25603) );
  NAND2_X1 U19074 ( .A1(n18338), .A2(n533), .ZN(n24451) );
  OAI22_X1 U19075 ( .A1(net716477), .A2(n24648), .B1(net767237), .B2(n548), 
        .ZN(n24459) );
  NAND2_X1 U19076 ( .A1(net767238), .A2(n24799), .ZN(n24468) );
  NAND2_X1 U19077 ( .A1(n18330), .A2(n531), .ZN(n24466) );
  AOI21_X1 U19078 ( .B1(net716417), .B2(n24762), .A(n24469), .ZN(n24464) );
  NAND2_X1 U19079 ( .A1(n18529), .A2(n528), .ZN(n24473) );
  OAI22_X1 U19080 ( .A1(n18316), .A2(n550), .B1(n551), .B2(n18315), .ZN(n24474) );
  NAND2_X1 U19081 ( .A1(net767239), .A2(n24722), .ZN(n24479) );
  AOI22_X1 U19082 ( .A1(n18307), .A2(n17712), .B1(net716405), .B2(n17711), 
        .ZN(n24478) );
  NAND2_X1 U19083 ( .A1(n18306), .A2(n538), .ZN(n24477) );
  NAND2_X1 U19084 ( .A1(n18311), .A2(n525), .ZN(n24481) );
  NAND2_X1 U19085 ( .A1(n18310), .A2(n539), .ZN(n24480) );
  INV_X1 U19086 ( .A(n25658), .ZN(n26678) );
  INV_X1 U19087 ( .A(n25612), .ZN(n26702) );
  AOI21_X1 U19088 ( .B1(n18300), .B2(n527), .A(n24463), .ZN(n24461) );
  AND2_X1 U19089 ( .A1(n25732), .A2(n25731), .ZN(n25649) );
  INV_X1 U19090 ( .A(n25666), .ZN(n26614) );
  AOI22_X1 U19091 ( .A1(n18330), .A2(n961), .B1(n18331), .B2(n17787), .ZN(
        n24503) );
  NAND2_X1 U19092 ( .A1(net767238), .A2(n24729), .ZN(n24502) );
  INV_X1 U19093 ( .A(n24083), .ZN(n24082) );
  AOI21_X1 U19094 ( .B1(n18300), .B2(n957), .A(n24510), .ZN(n24508) );
  NAND2_X1 U19095 ( .A1(n18529), .A2(n958), .ZN(n24515) );
  INV_X1 U19096 ( .A(n24073), .ZN(n24072) );
  OAI22_X1 U19097 ( .A1(n18316), .A2(n980), .B1(n981), .B2(n18315), .ZN(n24516) );
  AND2_X1 U19098 ( .A1(net767239), .A2(n24715), .ZN(n24522) );
  AOI22_X1 U19099 ( .A1(n18310), .A2(n969), .B1(n18311), .B2(n955), .ZN(n24520) );
  AND2_X1 U19100 ( .A1(net716405), .A2(n17789), .ZN(n24523) );
  OAI22_X1 U19101 ( .A1(net716477), .A2(n24641), .B1(net767237), .B2(n978), 
        .ZN(n24499) );
  NAND2_X1 U19102 ( .A1(n18338), .A2(n963), .ZN(n24491) );
  INV_X1 U19103 ( .A(n26441), .ZN(n26442) );
  AND2_X1 U19104 ( .A1(n25728), .A2(n25727), .ZN(n26753) );
  AND2_X1 U19105 ( .A1(n25730), .A2(n25729), .ZN(n26752) );
  AND2_X1 U19106 ( .A1(n25728), .A2(n25727), .ZN(n25645) );
  OR2_X1 U19107 ( .A1(n18332), .A2(n779), .ZN(n26277) );
  AND2_X1 U19108 ( .A1(n25728), .A2(n25727), .ZN(n25644) );
  NAND2_X1 U19109 ( .A1(n18339), .A2(n960), .ZN(n24494) );
  AND2_X1 U19110 ( .A1(n18347), .A2(n965), .ZN(n24495) );
  AND2_X1 U19111 ( .A1(n25693), .A2(n25692), .ZN(n25609) );
  AND2_X1 U19112 ( .A1(n25693), .A2(n25692), .ZN(n25608) );
  INV_X1 U19113 ( .A(net713726), .ZN(net713892) );
  AND2_X1 U19114 ( .A1(n25693), .A2(n25692), .ZN(n26772) );
  AND2_X1 U19115 ( .A1(n25707), .A2(n25706), .ZN(n26765) );
  AND2_X1 U19116 ( .A1(n18326), .A2(n24748), .ZN(n24506) );
  AND2_X1 U19117 ( .A1(n25707), .A2(n25706), .ZN(n25623) );
  AND2_X1 U19118 ( .A1(n25718), .A2(n25717), .ZN(n26758) );
  AND2_X1 U19119 ( .A1(net767235), .A2(n24749), .ZN(n24510) );
  AND2_X1 U19120 ( .A1(n25718), .A2(n25717), .ZN(n25634) );
  NAND2_X1 U19121 ( .A1(net716423), .A2(n17786), .ZN(n24507) );
  AND2_X1 U19122 ( .A1(n25718), .A2(n25717), .ZN(n25635) );
  AND2_X1 U19123 ( .A1(n18321), .A2(n966), .ZN(n24518) );
  NOR2_X1 U19124 ( .A1(net518461), .A2(n973), .ZN(n24517) );
  AND2_X1 U19125 ( .A1(n25743), .A2(n25742), .ZN(n25661) );
  AND2_X1 U19126 ( .A1(n25710), .A2(n25709), .ZN(n25626) );
  AND2_X1 U19127 ( .A1(n25743), .A2(n25742), .ZN(n25660) );
  AND2_X1 U19128 ( .A1(n25743), .A2(n25742), .ZN(n26745) );
  AND2_X1 U19129 ( .A1(n25710), .A2(n25709), .ZN(net717157) );
  AND2_X1 U19130 ( .A1(n25710), .A2(n25709), .ZN(n26763) );
  AND2_X1 U19131 ( .A1(n25730), .A2(n25729), .ZN(n25646) );
  AND2_X1 U19132 ( .A1(n25730), .A2(n25729), .ZN(n25647) );
  INV_X1 U19133 ( .A(n19338), .ZN(n25680) );
  INV_X1 U19134 ( .A(n26785), .ZN(n26609) );
  INV_X1 U19135 ( .A(n26776), .ZN(n18129) );
  AND2_X1 U19136 ( .A1(net715847), .A2(n25741), .ZN(n26746) );
  INV_X1 U19137 ( .A(net712961), .ZN(net709330) );
  AND2_X1 U19138 ( .A1(net715847), .A2(n25741), .ZN(n25658) );
  INV_X1 U19139 ( .A(n20042), .ZN(n26271) );
  AND2_X1 U19140 ( .A1(net715847), .A2(n25741), .ZN(n25659) );
  AND2_X1 U19141 ( .A1(n26776), .A2(n18166), .ZN(net741279) );
  NAND2_X1 U19142 ( .A1(n26776), .A2(net741565), .ZN(n26705) );
  AND2_X1 U19143 ( .A1(net715884), .A2(net715885), .ZN(n25629) );
  AND2_X1 U19144 ( .A1(net715884), .A2(net715885), .ZN(n26761) );
  INV_X1 U19145 ( .A(n24591), .ZN(n25675) );
  AND2_X1 U19146 ( .A1(n25712), .A2(n25711), .ZN(n26762) );
  INV_X1 U19147 ( .A(net518461), .ZN(net712520) );
  AND2_X1 U19148 ( .A1(n25736), .A2(n25735), .ZN(n26749) );
  OR2_X1 U19149 ( .A1(n18332), .A2(n897), .ZN(n24430) );
  OAI22_X1 U19150 ( .A1(n18362), .A2(n2084), .B1(n18361), .B2(n2085), .ZN(
        n24048) );
  AND2_X1 U19151 ( .A1(n25734), .A2(n25733), .ZN(n26750) );
  AND2_X1 U19152 ( .A1(n25712), .A2(n25711), .ZN(n25627) );
  AND2_X1 U19153 ( .A1(n25703), .A2(n25702), .ZN(n26767) );
  AND2_X1 U19154 ( .A1(n25734), .A2(n25733), .ZN(n25650) );
  AND2_X1 U19155 ( .A1(n25712), .A2(n25711), .ZN(n25628) );
  AND2_X1 U19156 ( .A1(n25734), .A2(n25733), .ZN(n25651) );
  AND2_X1 U19157 ( .A1(n25695), .A2(n25694), .ZN(n25611) );
  AND2_X1 U19158 ( .A1(n25697), .A2(n25696), .ZN(n26770) );
  AND2_X1 U19159 ( .A1(n25738), .A2(n25737), .ZN(n25655) );
  NAND2_X1 U19160 ( .A1(n18339), .A2(n530), .ZN(n24454) );
  INV_X1 U19161 ( .A(n24591), .ZN(n25676) );
  AND2_X1 U19162 ( .A1(n18347), .A2(n535), .ZN(n24455) );
  OAI22_X1 U19163 ( .A1(n18394), .A2(n2100), .B1(n2103), .B2(n18393), .ZN(
        n24058) );
  AND2_X1 U19164 ( .A1(n25720), .A2(n25719), .ZN(n26757) );
  AND2_X1 U19165 ( .A1(n25720), .A2(n25719), .ZN(n25636) );
  NOR2_X1 U19166 ( .A1(n18382), .A2(n2104), .ZN(n24057) );
  NAND2_X1 U19167 ( .A1(net767214), .A2(n17710), .ZN(n24462) );
  OAI22_X1 U19168 ( .A1(n18387), .A2(n2101), .B1(n24671), .B2(n18388), .ZN(
        n24060) );
  AND2_X1 U19169 ( .A1(net767235), .A2(n24763), .ZN(n24463) );
  OAI22_X1 U19170 ( .A1(n18318), .A2(n2082), .B1(n18390), .B2(n2097), .ZN(
        n24059) );
  NAND2_X1 U19171 ( .A1(net716423), .A2(n17708), .ZN(n24460) );
  AND2_X1 U19172 ( .A1(n25720), .A2(n25719), .ZN(n25637) );
  NAND2_X1 U19173 ( .A1(n18331), .A2(n17709), .ZN(n24467) );
  AND2_X1 U19174 ( .A1(n25703), .A2(n25702), .ZN(n25619) );
  AND2_X1 U19175 ( .A1(net767235), .A2(n17937), .ZN(n24061) );
  AND2_X1 U19176 ( .A1(n25703), .A2(n25702), .ZN(n25618) );
  AND2_X1 U19177 ( .A1(n25738), .A2(n25737), .ZN(n26748) );
  OR2_X1 U19178 ( .A1(n18332), .A2(n394), .ZN(n24439) );
  OR2_X1 U19179 ( .A1(n18332), .A2(n664), .ZN(n26655) );
  AND2_X1 U19180 ( .A1(n18321), .A2(n536), .ZN(n24483) );
  NOR2_X1 U19181 ( .A1(net518461), .A2(n543), .ZN(n24482) );
  AND2_X1 U19182 ( .A1(n25738), .A2(n25737), .ZN(n25654) );
  AND2_X1 U19183 ( .A1(n25701), .A2(n25700), .ZN(n25617) );
  AND2_X1 U19184 ( .A1(n25701), .A2(n25700), .ZN(n25616) );
  AND2_X1 U19185 ( .A1(n25701), .A2(n25700), .ZN(n26768) );
  OR2_X1 U19186 ( .A1(n18332), .A2(n703), .ZN(n26347) );
  AND2_X1 U19187 ( .A1(n25740), .A2(n25739), .ZN(n25657) );
  AND2_X1 U19188 ( .A1(n25740), .A2(n25739), .ZN(n25656) );
  AND2_X1 U19189 ( .A1(n25695), .A2(n25694), .ZN(n26771) );
  AND2_X1 U19190 ( .A1(n25716), .A2(n25715), .ZN(n26759) );
  AND2_X1 U19191 ( .A1(n25699), .A2(n25698), .ZN(n26769) );
  AND2_X1 U19192 ( .A1(n25716), .A2(n25715), .ZN(n25632) );
  AND2_X1 U19193 ( .A1(n25697), .A2(n25696), .ZN(n25613) );
  AND2_X1 U19194 ( .A1(n25716), .A2(n25715), .ZN(n25633) );
  AND2_X1 U19195 ( .A1(n25740), .A2(n25739), .ZN(n26747) );
  AND2_X1 U19196 ( .A1(n25697), .A2(n25696), .ZN(n25612) );
  AND2_X1 U19197 ( .A1(n25736), .A2(n25735), .ZN(n25652) );
  AND2_X1 U19198 ( .A1(n25699), .A2(n25698), .ZN(n25615) );
  INV_X1 U19199 ( .A(n18367), .ZN(net716491) );
  AND2_X1 U19200 ( .A1(n25699), .A2(n25698), .ZN(n25614) );
  AND2_X1 U19201 ( .A1(n25695), .A2(n25694), .ZN(n25610) );
  AND2_X1 U19202 ( .A1(n25736), .A2(n25735), .ZN(n25653) );
  INV_X1 U19203 ( .A(n19390), .ZN(n19308) );
  NOR3_X2 U19204 ( .A1(net366451), .A2(net366531), .A3(net716231), .ZN(
        net713863) );
  NAND2_X1 U19205 ( .A1(n18343), .A2(n524), .ZN(n24458) );
  OR2_X1 U19206 ( .A1(n19243), .A2(n19244), .ZN(net741541) );
  INV_X1 U19207 ( .A(n18158), .ZN(net720303) );
  OR2_X1 U19208 ( .A1(n20065), .A2(n20066), .ZN(n24614) );
  AND2_X1 U19209 ( .A1(n20076), .A2(n20060), .ZN(n24591) );
  OR2_X1 U19210 ( .A1(n20067), .A2(n20068), .ZN(n24615) );
  INV_X1 U19211 ( .A(n19385), .ZN(n19328) );
  INV_X1 U19212 ( .A(n19367), .ZN(n19337) );
  AND2_X1 U19213 ( .A1(n18325), .A2(n526), .ZN(n24469) );
  NOR2_X1 U19214 ( .A1(s_IFID_IR[28]), .A2(n25685), .ZN(n26776) );
  OR2_X1 U19215 ( .A1(n19245), .A2(n19246), .ZN(net741549) );
  AND2_X1 U19216 ( .A1(n20060), .A2(n20078), .ZN(n24619) );
  AND2_X1 U19217 ( .A1(n19255), .A2(n19238), .ZN(net741532) );
  NOR2_X1 U19218 ( .A1(n18395), .A2(n2106), .ZN(n24062) );
  NAND2_X1 U19219 ( .A1(n18343), .A2(n954), .ZN(n24498) );
  NOR2_X1 U19220 ( .A1(n26710), .A2(n6514), .ZN(n26709) );
  INV_X1 U19221 ( .A(n25662), .ZN(n26136) );
  NAND2_X1 U19222 ( .A1(n18329), .A2(n17788), .ZN(n24509) );
  AND2_X1 U19223 ( .A1(n19255), .A2(n19241), .ZN(net741539) );
  BUF_X2 U19224 ( .A(n19332), .Z(n24026) );
  INV_X1 U19225 ( .A(n19262), .ZN(net715842) );
  OR2_X1 U19226 ( .A1(n19248), .A2(n19249), .ZN(net741544) );
  INV_X1 U19227 ( .A(n19255), .ZN(net708964) );
  INV_X1 U19228 ( .A(net717087), .ZN(net767168) );
  AND2_X1 U19229 ( .A1(n20076), .A2(n20063), .ZN(n24617) );
  INV_X1 U19230 ( .A(n20117), .ZN(n25685) );
  OR2_X1 U19231 ( .A1(net716237), .A2(n1378), .ZN(n24832) );
  INV_X1 U19232 ( .A(n20049), .ZN(n26779) );
  INV_X1 U19233 ( .A(n20076), .ZN(n26778) );
  INV_X1 U19234 ( .A(n18138), .ZN(n25745) );
  INV_X1 U19235 ( .A(n20081), .ZN(n25744) );
  OR2_X1 U19236 ( .A1(n20069), .A2(n20070), .ZN(n24613) );
  AND2_X1 U19237 ( .A1(s_IFID_IR[27]), .A2(n19282), .ZN(n24813) );
  NOR2_X2 U19238 ( .A1(n24678), .A2(s_WB_MUX_CONTROL[1]), .ZN(net741608) );
  NOR2_X2 U19239 ( .A1(n24679), .A2(s_WB_MUX_CONTROL[0]), .ZN(n26663) );
  INV_X1 U19240 ( .A(net366479), .ZN(net716231) );
  NOR2_X1 U19241 ( .A1(n6746), .A2(n1498), .ZN(n26604) );
  OR2_X1 U19242 ( .A1(net787512), .A2(\core_inst/EXMEM_NPC/DFF_1/N3 ), .ZN(
        net740674) );
  NOR2_X2 U19243 ( .A1(n24679), .A2(s_WB_MUX_CONTROL[0]), .ZN(n25601) );
  NOR2_X2 U19244 ( .A1(s_WB_MUX_CONTROL[1]), .A2(s_WB_MUX_CONTROL[0]), .ZN(
        net741527) );
  NOR2_X2 U19245 ( .A1(n24678), .A2(s_WB_MUX_CONTROL[1]), .ZN(net741609) );
  AND2_X1 U19246 ( .A1(net366451), .A2(net366531), .ZN(net715584) );
  NOR2_X1 U19247 ( .A1(net750085), .A2(n4397), .ZN(n24027) );
  INV_X1 U19248 ( .A(n24028), .ZN(n24029) );
  BUF_X1 U19249 ( .A(n24028), .Z(n24305) );
  OAI22_X1 U19250 ( .A1(n24033), .A2(n23952), .B1(n26222), .B2(n24028), .ZN(
        net718103) );
  NAND3_X1 U19251 ( .A1(net716255), .A2(net717050), .A3(n26526), .ZN(n26527)
         );
  NAND3_X1 U19252 ( .A1(net716249), .A2(net712499), .A3(n26702), .ZN(n25545)
         );
  AND2_X1 U19253 ( .A1(net716255), .A2(n17956), .ZN(
        \core_inst/IDEX_NPC/DFF_5/N3 ) );
  NAND2_X1 U19254 ( .A1(n25853), .A2(n25854), .ZN(n26205) );
  NAND2_X1 U19255 ( .A1(n25851), .A2(n25850), .ZN(n26201) );
  XNOR2_X1 U19256 ( .A(n26205), .B(net716221), .ZN(n25979) );
  INV_X1 U19257 ( .A(net715048), .ZN(net766652) );
  NOR2_X1 U19258 ( .A1(n24266), .A2(net737907), .ZN(n26061) );
  OAI21_X1 U19259 ( .B1(n26728), .B2(net716263), .A(n26712), .ZN(n16384) );
  NAND2_X1 U19260 ( .A1(net749507), .A2(net749428), .ZN(net749476) );
  NAND2_X1 U19261 ( .A1(n25840), .A2(n24554), .ZN(n24031) );
  NOR2_X2 U19262 ( .A1(n24200), .A2(n24541), .ZN(n24557) );
  INV_X1 U19263 ( .A(n25622), .ZN(n26428) );
  AND2_X1 U19264 ( .A1(n25707), .A2(n25706), .ZN(n25622) );
  INV_X1 U19265 ( .A(net742576), .ZN(net765727) );
  AND2_X1 U19266 ( .A1(n25979), .A2(net713612), .ZN(n24032) );
  MUX2_X1 U19267 ( .A(n26098), .B(\core_inst/EXMEM_NPC/DFF_0/N3 ), .S(
        net741686), .Z(net755610) );
  NAND2_X1 U19268 ( .A1(n26235), .A2(net741603), .ZN(n26509) );
  XNOR2_X1 U19269 ( .A(n26208), .B(net716221), .ZN(n24191) );
  NOR2_X1 U19270 ( .A1(net714751), .A2(net718103), .ZN(n24034) );
  MUX2_X1 U19271 ( .A(n1182), .B(n26078), .S(net787528), .Z(n26180) );
  XNOR2_X1 U19272 ( .A(n25887), .B(net716215), .ZN(n24035) );
  BUF_X1 U19273 ( .A(net740075), .Z(net740076) );
  NAND2_X1 U19274 ( .A1(net741999), .A2(n24036), .ZN(n24486) );
  AND2_X1 U19275 ( .A1(net717052), .A2(n24487), .ZN(n24036) );
  INV_X1 U19276 ( .A(n25832), .ZN(n26210) );
  INV_X1 U19277 ( .A(net742576), .ZN(net765319) );
  MUX2_X2 U19278 ( .A(n26108), .B(\core_inst/EXMEM_NPC/DFF_2/N3 ), .S(
        net741686), .Z(net749725) );
  NAND2_X1 U19279 ( .A1(net715662), .A2(net750053), .ZN(n24037) );
  AOI21_X1 U19280 ( .B1(n24037), .B2(net740076), .A(net718033), .ZN(n24038) );
  AOI21_X1 U19281 ( .B1(n24037), .B2(net740076), .A(net718033), .ZN(net715647)
         );
  AOI21_X1 U19282 ( .B1(n24037), .B2(net740076), .A(net718033), .ZN(n24360) );
  NOR2_X1 U19283 ( .A1(net750085), .A2(n25339), .ZN(n25821) );
  XNOR2_X1 U19284 ( .A(n24039), .B(net716221), .ZN(n25828) );
  INV_X1 U19285 ( .A(net767320), .ZN(net749410) );
  NOR2_X1 U19286 ( .A1(n25503), .A2(net767320), .ZN(n26070) );
  NAND3_X1 U19287 ( .A1(net742368), .A2(net717048), .A3(n26490), .ZN(n24067)
         );
  AND2_X1 U19288 ( .A1(net742576), .A2(\core_inst/s_IF_OUT_IR_OUT [26]), .ZN(
        \core_inst/IFID_IR/DFF_26/N3 ) );
  OAI21_X1 U19289 ( .B1(net796114), .B2(n24066), .A(n24067), .ZN(
        \core_inst/IDEX_RF_IN1/DFF_1/N3 ) );
  OAI21_X1 U19290 ( .B1(net716333), .B2(n24076), .A(n24077), .ZN(
        \core_inst/IDEX_RF_IN1/DFF_11/N3 ) );
  NAND3_X1 U19291 ( .A1(n24054), .A2(n24055), .A3(n24056), .ZN(n24049) );
  NOR2_X1 U19292 ( .A1(net716369), .A2(n24041), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_6/N3 ) );
  NAND3_X1 U19293 ( .A1(n24065), .A2(n24529), .A3(n24283), .ZN(n26141) );
  AND2_X1 U19294 ( .A1(n24339), .A2(net733611), .ZN(n24065) );
  OAI22_X1 U19295 ( .A1(n19385), .A2(n2709), .B1(n26785), .B2(n25264), .ZN(
        n24073) );
  OAI22_X1 U19296 ( .A1(n19383), .A2(n2713), .B1(n19395), .B2(n2710), .ZN(
        n24074) );
  AOI21_X1 U19297 ( .B1(n19530), .B2(n24687), .A(n24074), .ZN(n24071) );
  NAND4_X1 U19298 ( .A1(n20021), .A2(n24075), .A3(n20022), .A4(n24070), .ZN(
        n24069) );
  NAND4_X1 U19299 ( .A1(n24071), .A2(n24072), .A3(n20031), .A4(n20036), .ZN(
        n24068) );
  OAI21_X1 U19300 ( .B1(n24068), .B2(n24069), .A(n26704), .ZN(n24066) );
  OAI22_X1 U19301 ( .A1(n19385), .A2(n3033), .B1(n26785), .B2(n25266), .ZN(
        n24083) );
  OAI22_X1 U19302 ( .A1(n19383), .A2(n3037), .B1(n19395), .B2(n3034), .ZN(
        n24084) );
  AOI21_X1 U19303 ( .B1(n19530), .B2(n24685), .A(n24084), .ZN(n24081) );
  NAND4_X1 U19304 ( .A1(n19979), .A2(n24085), .A3(n19980), .A4(n24080), .ZN(
        n24079) );
  NAND4_X1 U19305 ( .A1(n24081), .A2(n24082), .A3(n19989), .A4(n19994), .ZN(
        n24078) );
  OAI21_X1 U19306 ( .B1(n24078), .B2(n24079), .A(n26704), .ZN(n24076) );
  AND2_X1 U19307 ( .A1(net716257), .A2(n24263), .ZN(
        \core_inst/IFID_NPC/DFF_5/N3 ) );
  CLKBUF_X1 U19308 ( .A(net717830), .Z(net762759) );
  CLKBUF_X3 U19309 ( .A(net717060), .Z(net762754) );
  BUF_X1 U19310 ( .A(net713864), .Z(net717060) );
  AND2_X1 U19311 ( .A1(n25846), .A2(n26067), .ZN(n24086) );
  BUF_X1 U19312 ( .A(n26184), .Z(n24566) );
  CLKBUF_X1 U19313 ( .A(n26100), .Z(n24087) );
  BUF_X2 U19314 ( .A(net713560), .Z(net742507) );
  AND2_X1 U19315 ( .A1(net755033), .A2(n912), .ZN(n25440) );
  XNOR2_X1 U19316 ( .A(n26198), .B(net716215), .ZN(n24088) );
  CLKBUF_X1 U19317 ( .A(net715445), .Z(net755033) );
  OR2_X2 U19318 ( .A1(net714602), .A2(n25834), .ZN(n24089) );
  MUX2_X2 U19319 ( .A(n829), .B(n26105), .S(net787512), .Z(net749454) );
  OAI21_X1 U19320 ( .B1(net758037), .B2(n25972), .A(n24172), .ZN(n24090) );
  OAI21_X1 U19321 ( .B1(net758037), .B2(n25972), .A(n24172), .ZN(n24335) );
  INV_X1 U19322 ( .A(net713683), .ZN(net762660) );
  INV_X1 U19323 ( .A(net713683), .ZN(net762661) );
  CLKBUF_X1 U19324 ( .A(n23028), .Z(n24091) );
  OAI222_X1 U19325 ( .A1(n25599), .A2(n24277), .B1(n24310), .B2(net749387), 
        .C1(n24291), .C2(net762661), .ZN(n25915) );
  INV_X1 U19326 ( .A(net750182), .ZN(net762654) );
  BUF_X1 U19327 ( .A(n24570), .Z(n24098) );
  NOR2_X1 U19328 ( .A1(n25764), .A2(n25763), .ZN(n24092) );
  INV_X1 U19329 ( .A(n24265), .ZN(n24093) );
  MUX2_X2 U19330 ( .A(n24136), .B(n5585), .S(net741686), .Z(n24265) );
  NAND2_X1 U19331 ( .A1(n25514), .A2(n25578), .ZN(n24094) );
  BUF_X1 U19332 ( .A(n25995), .Z(n24552) );
  OAI222_X1 U19333 ( .A1(n26031), .A2(net749812), .B1(net762754), .B2(
        net749306), .C1(net717055), .C2(net749387), .ZN(n25879) );
  BUF_X1 U19334 ( .A(net718152), .Z(net762625) );
  CLKBUF_X1 U19335 ( .A(n24035), .Z(n24095) );
  CLKBUF_X1 U19336 ( .A(n26129), .Z(n24097) );
  OAI21_X1 U19337 ( .B1(n26129), .B2(n26128), .A(n26127), .ZN(net713811) );
  INV_X1 U19338 ( .A(net717543), .ZN(net762604) );
  INV_X1 U19339 ( .A(net755090), .ZN(net762597) );
  INV_X1 U19340 ( .A(n26732), .ZN(n24099) );
  NAND3_X1 U19343 ( .A1(net716249), .A2(n25665), .A3(n26648), .ZN(n24103) );
  AND2_X1 U19344 ( .A1(net716253), .A2(n13824), .ZN(
        \core_inst/IDEX_NPC/DFF_8/N3 ) );
  AND2_X1 U19345 ( .A1(net765341), .A2(n18055), .ZN(
        \core_inst/EXMEM_IR/DFF_12/N3 ) );
  NAND3_X1 U19346 ( .A1(net716261), .A2(net712397), .A3(n26600), .ZN(n26601)
         );
  OAI21_X1 U19347 ( .B1(net716377), .B2(n24102), .A(n24103), .ZN(
        \core_inst/IDEX_RF_IN1/DFF_15/N3 ) );
  OAI22_X1 U19348 ( .A1(n19385), .A2(n2889), .B1(n26785), .B2(n25268), .ZN(
        n24109) );
  OAI22_X1 U19349 ( .A1(n19383), .A2(n2893), .B1(n19395), .B2(n2890), .ZN(
        n24110) );
  AOI21_X1 U19350 ( .B1(n19530), .B2(n24689), .A(n24110), .ZN(n24107) );
  NAND4_X1 U19351 ( .A1(n19895), .A2(n24111), .A3(n19896), .A4(n24106), .ZN(
        n24105) );
  NAND4_X1 U19352 ( .A1(n24107), .A2(n24108), .A3(n19905), .A4(n19910), .ZN(
        n24104) );
  OAI21_X1 U19353 ( .B1(n24104), .B2(n24105), .A(n26704), .ZN(n24102) );
  NAND2_X1 U19354 ( .A1(net742017), .A2(n24587), .ZN(n25756) );
  NAND3_X1 U19355 ( .A1(n25754), .A2(n25753), .A3(n25756), .ZN(n25388) );
  NOR2_X1 U19356 ( .A1(n25755), .A2(n25388), .ZN(n26165) );
  OR2_X1 U19357 ( .A1(n25389), .A2(n22870), .ZN(n24329) );
  OR2_X2 U19358 ( .A1(n24329), .A2(net767203), .ZN(n25381) );
  NOR2_X1 U19359 ( .A1(net742243), .A2(net717087), .ZN(n24119) );
  MUX2_X1 U19360 ( .A(net713738), .B(net713726), .S(net742242), .Z(n24120) );
  OAI22_X1 U19361 ( .A1(n24338), .A2(net742271), .B1(n22949), .B2(n25663), 
        .ZN(n24121) );
  OAI22_X1 U19362 ( .A1(net717059), .A2(net767207), .B1(net717056), .B2(
        net748269), .ZN(n24122) );
  AND2_X1 U19363 ( .A1(n24269), .A2(n24119), .ZN(n24118) );
  NOR2_X1 U19364 ( .A1(n26219), .A2(net713728), .ZN(n24117) );
  NAND2_X1 U19365 ( .A1(n25381), .A2(n24120), .ZN(n24116) );
  OAI21_X1 U19366 ( .B1(n24121), .B2(n24122), .A(net713775), .ZN(n24114) );
  AOI211_X1 U19367 ( .C1(n24116), .C2(net750032), .A(n24117), .B(n24118), .ZN(
        n24115) );
  AND2_X1 U19368 ( .A1(n24115), .A2(n24114), .ZN(n24113) );
  NAND4_X1 U19369 ( .A1(n25776), .A2(n25775), .A3(n25774), .A4(n25773), .ZN(
        n24112) );
  OAI21_X1 U19370 ( .B1(n24112), .B2(net714182), .A(n24113), .ZN(n24399) );
  AND2_X1 U19371 ( .A1(net714494), .A2(n25999), .ZN(n26224) );
  INV_X1 U19372 ( .A(n26733), .ZN(n24123) );
  INV_X1 U19373 ( .A(n24326), .ZN(n26226) );
  INV_X1 U19374 ( .A(net716341), .ZN(net760161) );
  INV_X1 U19375 ( .A(net714585), .ZN(net760144) );
  BUF_X2 U19376 ( .A(n24175), .Z(n25579) );
  AOI21_X1 U19377 ( .B1(n25506), .B2(n25507), .A(net725577), .ZN(n24125) );
  AOI21_X1 U19378 ( .B1(n24235), .B2(net717091), .A(n24236), .ZN(n24126) );
  INV_X1 U19379 ( .A(n24258), .ZN(n24253) );
  INV_X1 U19381 ( .A(n24334), .ZN(n24128) );
  INV_X1 U19387 ( .A(n24126), .ZN(n24134) );
  NAND3_X1 U19388 ( .A1(\cu_inst/FW_UNIT/ITD_EXMEM/N17 ), .A2(n11743), .A3(
        n17659), .ZN(n24135) );
  AND2_X1 U19389 ( .A1(net742012), .A2(net715615), .ZN(net715443) );
  INV_X1 U19390 ( .A(net715445), .ZN(net742223) );
  INV_X1 U19391 ( .A(net715445), .ZN(net715420) );
  INV_X1 U19392 ( .A(net715445), .ZN(net718337) );
  NOR2_X1 U19393 ( .A1(net742223), .A2(n17859), .ZN(n25400) );
  OR2_X2 U19394 ( .A1(n24093), .A2(n24305), .ZN(n24138) );
  NAND2_X1 U19395 ( .A1(net750122), .A2(n25585), .ZN(n24137) );
  OR2_X1 U19396 ( .A1(n24137), .A2(net742241), .ZN(net717461) );
  BUF_X1 U19397 ( .A(n24137), .Z(n24140) );
  OR2_X1 U19398 ( .A1(n24137), .A2(net749697), .ZN(net755637) );
  OR2_X1 U19399 ( .A1(n24137), .A2(net749697), .ZN(net750277) );
  INV_X1 U19400 ( .A(net717461), .ZN(net749317) );
  NAND2_X1 U19401 ( .A1(net755258), .A2(net713733), .ZN(n25663) );
  AND3_X1 U19402 ( .A1(net753553), .A2(net714877), .A3(net714873), .ZN(
        net749427) );
  NAND3_X1 U19403 ( .A1(n25403), .A2(n25404), .A3(net755075), .ZN(net714354)
         );
  OAI22_X1 U19404 ( .A1(net714354), .A2(net714182), .B1(net714344), .B2(
        net714267), .ZN(n25970) );
  AND2_X1 U19405 ( .A1(net742275), .A2(n24333), .ZN(net728824) );
  OAI22_X1 U19406 ( .A1(net718361), .A2(net740717), .B1(net717105), .B2(n1696), 
        .ZN(n25387) );
  NAND2_X1 U19407 ( .A1(n23933), .A2(n24575), .ZN(net749841) );
  INV_X2 U19408 ( .A(n24140), .ZN(n26148) );
  AOI22_X1 U19409 ( .A1(n24544), .A2(n26148), .B1(net786856), .B2(net714249), 
        .ZN(n25900) );
  NAND3_X1 U19410 ( .A1(n24141), .A2(net714585), .A3(n25977), .ZN(n25982) );
  OR2_X1 U19411 ( .A1(n24528), .A2(net758037), .ZN(n24141) );
  OAI211_X1 U19412 ( .C1(net712872), .C2(n24089), .A(n24282), .B(n24335), .ZN(
        n24144) );
  OAI211_X1 U19413 ( .C1(net712872), .C2(n24089), .A(n24282), .B(n24090), .ZN(
        net755060) );
  NOR2_X1 U19414 ( .A1(n24144), .A2(net713964), .ZN(n24142) );
  NAND2_X1 U19415 ( .A1(net716261), .A2(s_IFID_IR[20]), .ZN(n26721) );
  INV_X1 U19416 ( .A(n26233), .ZN(n24143) );
  NAND2_X1 U19417 ( .A1(n26240), .A2(n24143), .ZN(n26235) );
  XNOR2_X1 U19418 ( .A(n26235), .B(net716223), .ZN(n26140) );
  NAND2_X1 U19419 ( .A1(n26140), .A2(n26405), .ZN(n26138) );
  NAND2_X1 U19420 ( .A1(net742368), .A2(s_IFID_IR[24]), .ZN(n26723) );
  NAND2_X1 U19421 ( .A1(net796255), .A2(s_IFID_IR[22]), .ZN(n26722) );
  OAI21_X1 U19422 ( .B1(n26723), .B2(n26705), .A(n24261), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_24/N3 ) );
  OAI21_X1 U19423 ( .B1(n26722), .B2(n26705), .A(n22874), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_22/N3 ) );
  NAND2_X1 U19424 ( .A1(n25447), .A2(n23896), .ZN(net714281) );
  NAND2_X1 U19425 ( .A1(net713467), .A2(net749442), .ZN(n25974) );
  NAND3_X1 U19426 ( .A1(n25980), .A2(net718380), .A3(n24571), .ZN(n24164) );
  NAND3_X1 U19427 ( .A1(n24164), .A2(net714585), .A3(n25981), .ZN(n24163) );
  NAND2_X1 U19428 ( .A1(n25991), .A2(net713892), .ZN(n24149) );
  NAND2_X1 U19429 ( .A1(n25990), .A2(net713736), .ZN(n24148) );
  OR2_X1 U19430 ( .A1(net749707), .A2(n24163), .ZN(n24165) );
  MUX2_X1 U19431 ( .A(n24148), .B(n24149), .S(net714559), .Z(n24147) );
  OAI22_X1 U19432 ( .A1(net755699), .A2(n24357), .B1(net796212), .B2(n25578), 
        .ZN(n24154) );
  OAI22_X1 U19433 ( .A1(net731327), .A2(net762754), .B1(net717055), .B2(
        net767206), .ZN(n24153) );
  OAI222_X1 U19434 ( .A1(n26031), .A2(net742259), .B1(n24303), .B2(net713773), 
        .C1(net750287), .C2(net713810), .ZN(n24152) );
  OR2_X1 U19435 ( .A1(n25471), .A2(n24425), .ZN(n24166) );
  INV_X1 U19436 ( .A(net713873), .ZN(net714575) );
  NAND2_X1 U19437 ( .A1(n25982), .A2(n24165), .ZN(n24162) );
  INV_X1 U19438 ( .A(net734346), .ZN(net755745) );
  OAI21_X1 U19439 ( .B1(n26229), .B2(net713738), .A(n24147), .ZN(n24146) );
  NOR2_X1 U19440 ( .A1(n26230), .A2(net713728), .ZN(n24145) );
  NOR3_X1 U19441 ( .A1(n24152), .A2(n24153), .A3(n24154), .ZN(n24151) );
  NAND2_X1 U19442 ( .A1(n24166), .A2(net732754), .ZN(n24150) );
  MUX2_X1 U19443 ( .A(net714401), .B(net713977), .S(net718367), .Z(n24157) );
  INV_X1 U19444 ( .A(n25921), .ZN(n24156) );
  MUX2_X1 U19445 ( .A(net714575), .B(n26000), .S(net718367), .Z(n24155) );
  NAND2_X1 U19446 ( .A1(net712872), .A2(net731199), .ZN(n24160) );
  NOR2_X1 U19447 ( .A1(n25978), .A2(n24327), .ZN(n24159) );
  NAND2_X1 U19448 ( .A1(n24162), .A2(n25984), .ZN(n24161) );
  NOR2_X1 U19449 ( .A1(n24327), .A2(n25978), .ZN(n24167) );
  AOI21_X1 U19450 ( .B1(n24150), .B2(n24151), .A(net713751), .ZN(net714553) );
  OAI22_X1 U19451 ( .A1(n24155), .A2(n24156), .B1(n24157), .B2(n24158), .ZN(
        net714552) );
  AOI21_X1 U19452 ( .B1(n24327), .B2(n25975), .A(net713154), .ZN(net725127) );
  NAND3_X1 U19453 ( .A1(n25974), .A2(n25975), .A3(net734346), .ZN(net725126)
         );
  AOI211_X1 U19454 ( .C1(n24160), .C2(net714585), .A(n25984), .B(net749542), 
        .ZN(net720370) );
  NAND2_X1 U19455 ( .A1(n24159), .A2(n25983), .ZN(net720368) );
  AOI21_X1 U19456 ( .B1(n24167), .B2(net755745), .A(n24161), .ZN(net720369) );
  CLKBUF_X1 U19457 ( .A(n24259), .Z(n24169) );
  BUF_X1 U19458 ( .A(net732533), .Z(net749274) );
  AND2_X1 U19459 ( .A1(net715170), .A2(net715169), .ZN(n24170) );
  AND2_X1 U19460 ( .A1(n22851), .A2(n24395), .ZN(n24171) );
  OR2_X1 U19461 ( .A1(net714559), .A2(n25833), .ZN(n24172) );
  CLKBUF_X1 U19462 ( .A(net713602), .Z(net755740) );
  INV_X1 U19463 ( .A(net713777), .ZN(net713602) );
  INV_X1 U19464 ( .A(n24179), .ZN(n25871) );
  OAI21_X1 U19465 ( .B1(n25366), .B2(n26130), .A(n24096), .ZN(net755714) );
  INV_X1 U19466 ( .A(net716341), .ZN(net755708) );
  CLKBUF_X1 U19467 ( .A(n25861), .Z(n24173) );
  INV_X1 U19468 ( .A(n26175), .ZN(n26176) );
  OR3_X1 U19469 ( .A1(n26241), .A2(n25395), .A3(n25396), .ZN(n24542) );
  INV_X1 U19470 ( .A(n25781), .ZN(n25785) );
  AND2_X1 U19471 ( .A1(net718372), .A2(net750182), .ZN(n24176) );
  NAND2_X1 U19472 ( .A1(n25899), .A2(n25900), .ZN(n24177) );
  OR2_X2 U19473 ( .A1(n24276), .A2(net796258), .ZN(n24560) );
  OR2_X2 U19474 ( .A1(net714689), .A2(net750255), .ZN(n24276) );
  INV_X1 U19475 ( .A(net713561), .ZN(net713606) );
  XNOR2_X1 U19476 ( .A(n26052), .B(net366479), .ZN(n24179) );
  OAI21_X1 U19487 ( .B1(n26118), .B2(n24354), .A(n24557), .ZN(net749338) );
  INV_X1 U19488 ( .A(n24557), .ZN(n24562) );
  AOI22_X1 U19489 ( .A1(net714249), .A2(n24277), .B1(net750057), .B2(net742157), .ZN(n25451) );
  INV_X1 U19490 ( .A(net718086), .ZN(net718087) );
  NAND2_X1 U19491 ( .A1(n25419), .A2(net742092), .ZN(n25421) );
  NOR2_X1 U19492 ( .A1(n24271), .A2(net767203), .ZN(n25921) );
  OAI222_X1 U19493 ( .A1(n24560), .A2(net755238), .B1(net750287), .B2(
        net749525), .C1(n24291), .C2(net748269), .ZN(n25881) );
  INV_X1 U19494 ( .A(n25780), .ZN(n24190) );
  INV_X1 U19495 ( .A(n25780), .ZN(n25788) );
  MUX2_X1 U19496 ( .A(\core_inst/EXMEM_NPC/DFF_4/N3 ), .B(n26096), .S(
        net787528), .Z(net713687) );
  INV_X1 U19497 ( .A(net749465), .ZN(net755260) );
  INV_X1 U19498 ( .A(net755637), .ZN(net755258) );
  INV_X1 U19499 ( .A(net714559), .ZN(net755241) );
  INV_X1 U19500 ( .A(net714559), .ZN(net755240) );
  BUF_X1 U19501 ( .A(n24575), .Z(n24277) );
  BUF_X1 U19502 ( .A(n26184), .Z(n24567) );
  NOR2_X1 U19503 ( .A1(net715551), .A2(n25469), .ZN(n24194) );
  BUF_X1 U19504 ( .A(net750024), .Z(net749967) );
  CLKBUF_X1 U19505 ( .A(n26098), .Z(n24195) );
  OAI22_X1 U19506 ( .A1(n26080), .A2(net741686), .B1(net716237), .B2(
        \core_inst/EXMEM_NPC/DFF_27/N3 ), .ZN(net755216) );
  AND2_X2 U19507 ( .A1(net737672), .A2(net715632), .ZN(n25390) );
  NOR2_X1 U19508 ( .A1(n26035), .A2(net713669), .ZN(net755210) );
  BUF_X1 U19509 ( .A(net749698), .Z(net755207) );
  AND2_X1 U19510 ( .A1(n25587), .A2(n24576), .ZN(n24346) );
  BUF_X1 U19511 ( .A(net749338), .Z(net755137) );
  INV_X1 U19512 ( .A(n24525), .ZN(n24196) );
  BUF_X1 U19513 ( .A(n23970), .Z(n25586) );
  INV_X1 U19514 ( .A(n25941), .ZN(n25980) );
  INV_X1 U19515 ( .A(n25586), .ZN(n24422) );
  NAND2_X1 U19516 ( .A1(n25586), .A2(n24420), .ZN(n24419) );
  INV_X1 U19517 ( .A(n24199), .ZN(n24198) );
  INV_X1 U19518 ( .A(net749410), .ZN(net755086) );
  AND2_X1 U19519 ( .A1(n25979), .A2(net713612), .ZN(n24200) );
  BUF_X1 U19520 ( .A(net737672), .Z(net749951) );
  NAND2_X1 U19521 ( .A1(n25851), .A2(n25850), .ZN(n24201) );
  INV_X1 U19522 ( .A(net713990), .ZN(net755056) );
  CLKBUF_X1 U19523 ( .A(net713740), .Z(net755048) );
  AND2_X1 U19524 ( .A1(n24178), .A2(n24274), .ZN(n24202) );
  BUF_X2 U19525 ( .A(net713636), .Z(net742315) );
  BUF_X2 U19526 ( .A(net762625), .Z(net750255) );
  AND2_X1 U19527 ( .A1(net755056), .A2(net715284), .ZN(n24203) );
  OAI222_X1 U19528 ( .A1(n24310), .A2(net755238), .B1(net713851), .B2(n24269), 
        .C1(net713907), .C2(net742271), .ZN(n26030) );
  AND2_X1 U19529 ( .A1(n25854), .A2(n22667), .ZN(n24204) );
  NOR2_X1 U19530 ( .A1(n25746), .A2(n25370), .ZN(net717926) );
  INV_X1 U19531 ( .A(n25589), .ZN(n25590) );
  OR2_X1 U19532 ( .A1(n25885), .A2(n24205), .ZN(n25891) );
  OR2_X1 U19533 ( .A1(n25886), .A2(net767210), .ZN(n24205) );
  OR2_X1 U19534 ( .A1(net780522), .A2(n25384), .ZN(n24206) );
  CLKBUF_X1 U19535 ( .A(net731713), .Z(net754997) );
  CLKBUF_X1 U19536 ( .A(n26132), .Z(n24292) );
  INV_X1 U19537 ( .A(net712365), .ZN(net754762) );
  INV_X1 U19539 ( .A(n26729), .ZN(n24209) );
  INV_X1 U19540 ( .A(n24787), .ZN(n24210) );
  INV_X1 U19541 ( .A(n26737), .ZN(n24211) );
  INV_X1 U19542 ( .A(n26735), .ZN(n24212) );
  INV_X1 U19543 ( .A(net718082), .ZN(net718083) );
  CLKBUF_X1 U19544 ( .A(net718083), .Z(net749817) );
  NOR2_X1 U19545 ( .A1(net714751), .A2(net718103), .ZN(net739130) );
  NAND2_X1 U19546 ( .A1(net755214), .A2(net762625), .ZN(n25418) );
  NOR2_X1 U19547 ( .A1(net728314), .A2(net742324), .ZN(n24228) );
  OAI22_X1 U19548 ( .A1(net717056), .A2(net717875), .B1(net713907), .B2(
        net750274), .ZN(n24230) );
  OAI22_X1 U19549 ( .A1(net717053), .A2(net750093), .B1(net785219), .B2(
        net755238), .ZN(n24229) );
  OAI22_X1 U19550 ( .A1(n24310), .A2(n24277), .B1(n26031), .B2(n24577), .ZN(
        n24231) );
  OAI222_X1 U19551 ( .A1(net742483), .A2(n24233), .B1(n25443), .B2(net762661), 
        .C1(net713753), .C2(net717059), .ZN(n24225) );
  NOR2_X1 U19552 ( .A1(n24291), .A2(net749260), .ZN(n24224) );
  NOR3_X1 U19553 ( .A1(n24229), .A2(n24230), .A3(n24228), .ZN(n24227) );
  INV_X1 U19554 ( .A(n24231), .ZN(n24226) );
  NOR2_X1 U19555 ( .A1(n24224), .A2(n24225), .ZN(n24223) );
  NAND2_X1 U19556 ( .A1(n24570), .A2(net736366), .ZN(n24222) );
  NAND2_X1 U19557 ( .A1(n26054), .A2(net739078), .ZN(n24219) );
  NOR2_X1 U19558 ( .A1(n25994), .A2(net713726), .ZN(n24216) );
  NOR2_X1 U19559 ( .A1(n24565), .A2(net717087), .ZN(n24215) );
  OAI211_X1 U19560 ( .C1(n26063), .C2(net748269), .A(n24226), .B(n24227), .ZN(
        n24220) );
  OAI211_X1 U19561 ( .C1(n24539), .C2(net717074), .A(n24222), .B(n24223), .ZN(
        n24221) );
  NOR2_X1 U19562 ( .A1(n25579), .A2(net713751), .ZN(n24218) );
  OAI21_X1 U19563 ( .B1(n25374), .B2(net739078), .A(n24219), .ZN(n24217) );
  OAI22_X1 U19564 ( .A1(net713728), .A2(n26191), .B1(n26192), .B2(n25662), 
        .ZN(n24214) );
  MUX2_X1 U19565 ( .A(n24215), .B(n24216), .S(n24547), .Z(n24213) );
  AND3_X1 U19566 ( .A1(net755075), .A2(n25404), .A3(n25403), .ZN(n24232) );
  OAI21_X1 U19567 ( .B1(n24221), .B2(n24220), .A(net713775), .ZN(net746315) );
  OAI21_X1 U19568 ( .B1(n24217), .B2(n26059), .A(n24218), .ZN(net714506) );
  NAND2_X1 U19569 ( .A1(n26028), .A2(net767208), .ZN(net714508) );
  AOI211_X1 U19570 ( .C1(n24232), .C2(net714306), .A(n24213), .B(n24214), .ZN(
        net714507) );
  NOR2_X1 U19571 ( .A1(n26040), .A2(net749709), .ZN(n24234) );
  OR2_X1 U19572 ( .A1(n26040), .A2(net767209), .ZN(n24238) );
  OAI22_X1 U19573 ( .A1(n25595), .A2(n4343), .B1(net738474), .B2(n24815), .ZN(
        net715528) );
  NAND2_X1 U19574 ( .A1(n25585), .A2(net718152), .ZN(n25782) );
  NOR2_X1 U19575 ( .A1(n25782), .A2(net717511), .ZN(net731344) );
  NAND2_X1 U19576 ( .A1(net750025), .A2(net749454), .ZN(n25770) );
  MUX2_X1 U19577 ( .A(net767234), .B(net713736), .S(n26188), .Z(n24251) );
  INV_X1 U19578 ( .A(net749822), .ZN(net736366) );
  MUX2_X1 U19579 ( .A(net713892), .B(n26136), .S(n26188), .Z(n24252) );
  NOR2_X1 U19580 ( .A1(net728314), .A2(net742483), .ZN(n24257) );
  OAI22_X1 U19581 ( .A1(net717075), .A2(n24269), .B1(net717055), .B2(net762661), .ZN(n24256) );
  OAI22_X1 U19582 ( .A1(n24310), .A2(net748269), .B1(net762753), .B2(net755238), .ZN(n24258) );
  NAND2_X1 U19583 ( .A1(net714309), .A2(n25858), .ZN(n24244) );
  NAND3_X1 U19584 ( .A1(n25857), .A2(net715027), .A3(n25856), .ZN(n24243) );
  INV_X1 U19585 ( .A(net715018), .ZN(net736356) );
  NAND2_X1 U19586 ( .A1(net749822), .A2(n24251), .ZN(n24250) );
  OAI21_X1 U19587 ( .B1(n26038), .B2(n24252), .A(net736366), .ZN(n24249) );
  NAND2_X1 U19588 ( .A1(net712466), .A2(n24359), .ZN(n24255) );
  NOR2_X1 U19589 ( .A1(n24256), .A2(n24257), .ZN(n24254) );
  NOR4_X1 U19590 ( .A1(n25859), .A2(n24243), .A3(n24244), .A4(n24245), .ZN(
        n24242) );
  NOR4_X1 U19591 ( .A1(net714182), .A2(net715015), .A3(net736356), .A4(n24246), 
        .ZN(n24241) );
  NAND2_X1 U19592 ( .A1(n24249), .A2(n24250), .ZN(n24248) );
  NAND3_X1 U19593 ( .A1(n24253), .A2(n24254), .A3(n24255), .ZN(n24247) );
  AOI21_X1 U19594 ( .B1(n24241), .B2(net749839), .A(n24242), .ZN(n24240) );
  NAND2_X1 U19595 ( .A1(n24545), .A2(net767208), .ZN(n24237) );
  AOI21_X1 U19596 ( .B1(n24247), .B2(net713775), .A(n24248), .ZN(n24239) );
  NAND4_X1 U19597 ( .A1(n24239), .A2(n24238), .A3(n24237), .A4(n24240), .ZN(
        n24236) );
  OR2_X1 U19598 ( .A1(n24570), .A2(net749500), .ZN(n24425) );
  NAND2_X1 U19599 ( .A1(net749500), .A2(n24311), .ZN(n25860) );
  NAND2_X1 U19600 ( .A1(net749500), .A2(net749454), .ZN(n26158) );
  NAND2_X1 U19601 ( .A1(n26120), .A2(net749902), .ZN(net712855) );
  AND4_X1 U19602 ( .A1(n24169), .A2(n25762), .A3(n25774), .A4(n25761), .ZN(
        n25596) );
  NAND4_X1 U19603 ( .A1(n24259), .A2(n25762), .A3(n25774), .A4(n25761), .ZN(
        n24342) );
  INV_X1 U19604 ( .A(net742612), .ZN(net716353) );
  NAND2_X1 U19605 ( .A1(n24261), .A2(n24535), .ZN(n6695) );
  OAI21_X1 U19606 ( .B1(n26720), .B2(n26705), .A(n22874), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_16/N3 ) );
  OAI21_X1 U19607 ( .B1(n26569), .B2(n26705), .A(n24261), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_17/N3 ) );
  OAI21_X1 U19608 ( .B1(n26577), .B2(n26705), .A(n24261), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_19/N3 ) );
  OAI21_X1 U19609 ( .B1(n26721), .B2(n26705), .A(n22874), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_20/N3 ) );
  OAI21_X1 U19610 ( .B1(net712384), .B2(n26705), .A(n22874), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_21/N3 ) );
  NAND2_X1 U19611 ( .A1(n24261), .A2(n24535), .ZN(n24573) );
  AOI21_X1 U19612 ( .B1(n6514), .B2(n26710), .A(n26709), .ZN(n24263) );
  INV_X1 U19613 ( .A(n26201), .ZN(n26199) );
  INV_X1 U19614 ( .A(n25991), .ZN(n25990) );
  CLKBUF_X1 U19615 ( .A(n25392), .Z(n24264) );
  AND2_X1 U19616 ( .A1(n25444), .A2(n25445), .ZN(n26009) );
  CLKBUF_X3 U19617 ( .A(net712893), .Z(net750287) );
  OR2_X1 U19618 ( .A1(net717543), .A2(net755207), .ZN(n24266) );
  NAND2_X1 U19619 ( .A1(n26090), .A2(net716237), .ZN(n24268) );
  INV_X1 U19620 ( .A(n24192), .ZN(n24269) );
  INV_X1 U19621 ( .A(n25381), .ZN(n26038) );
  INV_X1 U19622 ( .A(net715359), .ZN(net750264) );
  OAI222_X1 U19623 ( .A1(net717055), .A2(n24277), .B1(n24546), .B2(net748269), 
        .C1(n24233), .C2(n24358), .ZN(n26033) );
  NOR2_X1 U19624 ( .A1(net765428), .A2(net742243), .ZN(n24272) );
  CLKBUF_X3 U19625 ( .A(net713612), .Z(net750238) );
  AOI21_X1 U19626 ( .B1(n25939), .B2(net742423), .A(n25373), .ZN(n24273) );
  MUX2_X1 U19627 ( .A(net742224), .B(n367), .S(net741686), .Z(net750228) );
  NAND2_X2 U19628 ( .A1(n25367), .A2(n24832), .ZN(n24274) );
  AND2_X1 U19629 ( .A1(net737672), .A2(net715632), .ZN(n24275) );
  NAND2_X1 U19630 ( .A1(n25367), .A2(n24832), .ZN(net713669) );
  AND2_X1 U19631 ( .A1(net737672), .A2(net715632), .ZN(net742284) );
  INV_X1 U19632 ( .A(n26208), .ZN(n26076) );
  MUX2_X1 U19633 ( .A(n25392), .B(n17924), .S(net741686), .Z(n24575) );
  INV_X1 U19634 ( .A(n26047), .ZN(n25429) );
  OR2_X1 U19635 ( .A1(net749273), .A2(net742243), .ZN(net750203) );
  INV_X1 U19636 ( .A(n24265), .ZN(n24279) );
  INV_X1 U19637 ( .A(n24265), .ZN(n24278) );
  XNOR2_X1 U19638 ( .A(n24312), .B(net716215), .ZN(n24299) );
  AND2_X2 U19639 ( .A1(n25839), .A2(n25838), .ZN(n24312) );
  OR2_X1 U19640 ( .A1(net718351), .A2(n5618), .ZN(n25386) );
  CLKBUF_X1 U19641 ( .A(net717510), .Z(net750176) );
  NAND2_X1 U19642 ( .A1(n25515), .A2(n25993), .ZN(n24282) );
  NAND2_X1 U19643 ( .A1(n24543), .A2(n25442), .ZN(n26019) );
  AND2_X2 U19644 ( .A1(net747347), .A2(net747343), .ZN(net750158) );
  AND2_X1 U19645 ( .A1(net747347), .A2(net747343), .ZN(n24401) );
  BUF_X1 U19646 ( .A(n24034), .Z(n24283) );
  INV_X1 U19647 ( .A(n26000), .ZN(n26137) );
  INV_X1 U19648 ( .A(n23979), .ZN(n24286) );
  CLKBUF_X1 U19649 ( .A(n24551), .Z(n24287) );
  INV_X1 U19650 ( .A(net717543), .ZN(net714249) );
  CLKBUF_X1 U19651 ( .A(n22873), .Z(n24289) );
  OR2_X1 U19652 ( .A1(n25823), .A2(n25898), .ZN(n24290) );
  AOI21_X1 U19653 ( .B1(n25506), .B2(n25507), .A(net725577), .ZN(n25505) );
  INV_X1 U19654 ( .A(net731329), .ZN(net750090) );
  INV_X1 U19655 ( .A(net713894), .ZN(net713978) );
  BUF_X1 U19656 ( .A(net713560), .Z(net742506) );
  INV_X1 U19657 ( .A(n24204), .ZN(n24293) );
  CLKBUF_X1 U19658 ( .A(n25393), .Z(n24294) );
  BUF_X2 U19659 ( .A(n24569), .Z(n24295) );
  XNOR2_X1 U19660 ( .A(n24201), .B(net716221), .ZN(n24296) );
  NOR3_X2 U19661 ( .A1(n25870), .A2(n25869), .A3(n25868), .ZN(n26724) );
  OR2_X1 U19662 ( .A1(net755060), .A2(net713964), .ZN(n24297) );
  AOI21_X1 U19663 ( .B1(net742011), .B2(net780579), .A(net717926), .ZN(
        net718092) );
  NOR2_X1 U19664 ( .A1(n24323), .A2(n25505), .ZN(n24298) );
  INV_X1 U19665 ( .A(net750274), .ZN(net750032) );
  BUF_X1 U19666 ( .A(net731344), .Z(net750025) );
  INV_X1 U19667 ( .A(net717845), .ZN(net717510) );
  INV_X1 U19668 ( .A(net713882), .ZN(net713779) );
  CLKBUF_X1 U19669 ( .A(n26172), .Z(n24355) );
  NAND2_X1 U19670 ( .A1(n25921), .A2(n24294), .ZN(net713897) );
  INV_X1 U19671 ( .A(n26052), .ZN(n26051) );
  XNOR2_X1 U19672 ( .A(\cu_inst/FW_UNIT/ITD_EXMEM/N17 ), .B(n24574), .ZN(
        net715769) );
  CLKBUF_X1 U19673 ( .A(net749317), .Z(net749898) );
  AOI21_X1 U19674 ( .B1(n26110), .B2(net716237), .A(n25470), .ZN(net749993) );
  AOI21_X1 U19675 ( .B1(n24194), .B2(net716237), .A(n25470), .ZN(n24301) );
  AOI21_X1 U19676 ( .B1(n26110), .B2(net716237), .A(n25470), .ZN(n26193) );
  BUF_X1 U19677 ( .A(net715794), .Z(net749987) );
  NOR2_X1 U19678 ( .A1(\cu_inst/FW_UNIT/ITD_EXMEM/N17 ), .A2(
        \cu_inst/FW_UNIT/ITD_EXMEM/N14 ), .ZN(net715794) );
  INV_X1 U19679 ( .A(n22845), .ZN(n25945) );
  INV_X1 U19680 ( .A(net717056), .ZN(net712468) );
  NAND2_X1 U19681 ( .A1(n25921), .A2(net718367), .ZN(net749977) );
  CLKBUF_X3 U19682 ( .A(net717103), .Z(net749972) );
  CLKBUF_X3 U19683 ( .A(n24377), .Z(n24303) );
  INV_X1 U19684 ( .A(net713810), .ZN(net749936) );
  INV_X2 U19685 ( .A(net713151), .ZN(net713810) );
  AND2_X1 U19686 ( .A1(n24269), .A2(net742243), .ZN(n24304) );
  BUF_X1 U19687 ( .A(net714977), .Z(net749930) );
  NOR2_X2 U19688 ( .A1(net718349), .A2(n26168), .ZN(n26233) );
  INV_X1 U19689 ( .A(net742339), .ZN(net749910) );
  AND2_X1 U19690 ( .A1(n25784), .A2(n25783), .ZN(n24306) );
  NAND2_X1 U19691 ( .A1(n25942), .A2(n25981), .ZN(net749905) );
  OR2_X1 U19692 ( .A1(n24403), .A2(n26068), .ZN(n24307) );
  CLKBUF_X3 U19693 ( .A(n24377), .Z(n24310) );
  OR2_X1 U19694 ( .A1(n24192), .A2(n23977), .ZN(n24308) );
  MUX2_X2 U19695 ( .A(n26085), .B(\core_inst/EXMEM_NPC/DFF_30/N3 ), .S(
        net741686), .Z(net713151) );
  NAND2_X1 U19696 ( .A1(net780598), .A2(net740674), .ZN(n24358) );
  CLKBUF_X1 U19697 ( .A(net717543), .Z(net742304) );
  OAI222_X1 U19698 ( .A1(net750287), .A2(net749823), .B1(net717074), .B2(
        net717875), .C1(net755757), .C2(net749387), .ZN(n26029) );
  INV_X1 U19699 ( .A(n24279), .ZN(n24311) );
  INV_X1 U19700 ( .A(n26222), .ZN(n24544) );
  AND2_X1 U19701 ( .A1(net713707), .A2(n24285), .ZN(n26183) );
  INV_X1 U19702 ( .A(net786844), .ZN(net749832) );
  INV_X1 U19703 ( .A(net713672), .ZN(net749820) );
  INV_X1 U19704 ( .A(net749820), .ZN(net749822) );
  OR2_X1 U19705 ( .A1(n24095), .A2(n24301), .ZN(n24313) );
  OR2_X1 U19706 ( .A1(n24035), .A2(net749993), .ZN(net749798) );
  NAND2_X1 U19707 ( .A1(net749372), .A2(net713740), .ZN(n26134) );
  INV_X1 U19708 ( .A(n23972), .ZN(n26188) );
  INV_X1 U19709 ( .A(n24574), .ZN(n24316) );
  INV_X1 U19710 ( .A(net767357), .ZN(net713672) );
  OAI21_X1 U19711 ( .B1(n24346), .B2(n26041), .A(n24197), .ZN(n24317) );
  INV_X1 U19712 ( .A(net713681), .ZN(net749732) );
  INV_X1 U19713 ( .A(net715032), .ZN(net715200) );
  AND2_X1 U19714 ( .A1(n25822), .A2(n23976), .ZN(n24318) );
  INV_X1 U19715 ( .A(net714309), .ZN(net749709) );
  INV_X1 U19716 ( .A(net749709), .ZN(net749710) );
  NAND2_X1 U19717 ( .A1(n24528), .A2(n25943), .ZN(n24319) );
  NAND2_X1 U19718 ( .A1(n24528), .A2(n25943), .ZN(net749707) );
  INV_X1 U19719 ( .A(n23967), .ZN(n26194) );
  INV_X1 U19720 ( .A(net713867), .ZN(net749685) );
  INV_X1 U19721 ( .A(net750158), .ZN(net749679) );
  INV_X1 U19722 ( .A(net749369), .ZN(net749664) );
  INV_X1 U19723 ( .A(net742284), .ZN(net742209) );
  NOR2_X1 U19724 ( .A1(net717510), .A2(n25782), .ZN(n24321) );
  AND3_X1 U19725 ( .A1(net742092), .A2(n26143), .A3(n24206), .ZN(n24322) );
  NAND3_X1 U19726 ( .A1(n25508), .A2(n25416), .A3(n23822), .ZN(n24323) );
  MUX2_X2 U19727 ( .A(n26106), .B(\core_inst/EXMEM_NPC/DFF_28/N3 ), .S(
        net741686), .Z(net713564) );
  AND2_X1 U19728 ( .A1(net762654), .A2(net749832), .ZN(n24324) );
  CLKBUF_X1 U19729 ( .A(n26101), .Z(n24325) );
  XNOR2_X1 U19730 ( .A(n23028), .B(net716223), .ZN(net749636) );
  NAND2_X1 U19731 ( .A1(net755216), .A2(n24552), .ZN(n24326) );
  INV_X1 U19732 ( .A(net755216), .ZN(net714494) );
  INV_X1 U19733 ( .A(n25873), .ZN(n26128) );
  NOR2_X1 U19734 ( .A1(n25438), .A2(net728159), .ZN(n24327) );
  INV_X1 U19735 ( .A(net713554), .ZN(net713967) );
  AND2_X1 U19736 ( .A1(n24178), .A2(n24274), .ZN(net714861) );
  INV_X1 U19737 ( .A(net713669), .ZN(net714251) );
  OR2_X1 U19738 ( .A1(n25791), .A2(n25792), .ZN(n24328) );
  OR3_X1 U19739 ( .A1(net716341), .A2(n24610), .A3(n26705), .ZN(n24535) );
  MUX2_X2 U19740 ( .A(n26108), .B(\core_inst/EXMEM_NPC/DFF_2/N3 ), .S(
        net741686), .Z(net713683) );
  INV_X1 U19741 ( .A(n24195), .ZN(n26102) );
  NAND2_X1 U19742 ( .A1(n25425), .A2(n25426), .ZN(n24330) );
  NAND2_X1 U19743 ( .A1(net713923), .A2(n25993), .ZN(n26561) );
  CLKBUF_X1 U19744 ( .A(n25447), .Z(n24332) );
  AND2_X1 U19745 ( .A1(net749841), .A2(net715032), .ZN(n24333) );
  CLKBUF_X1 U19746 ( .A(net742242), .Z(net749534) );
  NAND2_X1 U19747 ( .A1(n26073), .A2(net713813), .ZN(net749533) );
  AND2_X1 U19748 ( .A1(net738443), .A2(net713833), .ZN(net717547) );
  NAND2_X1 U19749 ( .A1(net749489), .A2(net713740), .ZN(n24338) );
  INV_X1 U19750 ( .A(n26186), .ZN(n26189) );
  AND2_X1 U19751 ( .A1(net714559), .A2(n25833), .ZN(n25972) );
  INV_X1 U19752 ( .A(net714559), .ZN(net713906) );
  INV_X1 U19753 ( .A(net755637), .ZN(net749489) );
  INV_X1 U19754 ( .A(net749542), .ZN(net714603) );
  CLKBUF_X1 U19755 ( .A(n23029), .Z(n24340) );
  NAND2_X1 U19756 ( .A1(net755214), .A2(net742242), .ZN(net749465) );
  NOR2_X1 U19757 ( .A1(n25389), .A2(n22870), .ZN(net737713) );
  INV_X1 U19758 ( .A(net742265), .ZN(net749443) );
  NOR2_X1 U19759 ( .A1(n26459), .A2(n5577), .ZN(n26574) );
  INV_X1 U19760 ( .A(n26190), .ZN(n26213) );
  AND2_X1 U19761 ( .A1(net718349), .A2(n26168), .ZN(n26234) );
  INV_X1 U19762 ( .A(n26096), .ZN(n26097) );
  AND2_X1 U19763 ( .A1(net737713), .A2(net713773), .ZN(n25380) );
  NOR2_X1 U19764 ( .A1(n24270), .A2(net713773), .ZN(n24411) );
  INV_X1 U19765 ( .A(net714476), .ZN(net732754) );
  INV_X1 U19766 ( .A(net713773), .ZN(net734022) );
  AND2_X1 U19767 ( .A1(n24345), .A2(n25852), .ZN(n24344) );
  NAND2_X1 U19768 ( .A1(n24268), .A2(n24608), .ZN(n24345) );
  XNOR2_X1 U19769 ( .A(n26181), .B(net716223), .ZN(n24347) );
  INV_X1 U19770 ( .A(n26132), .ZN(n24348) );
  INV_X1 U19771 ( .A(net767357), .ZN(net731329) );
  BUF_X1 U19772 ( .A(n26065), .Z(n24576) );
  OR2_X1 U19773 ( .A1(net713829), .A2(net713151), .ZN(n24830) );
  INV_X1 U19774 ( .A(net713151), .ZN(net748274) );
  INV_X1 U19775 ( .A(n26197), .ZN(n26200) );
  OR2_X1 U19776 ( .A1(n24571), .A2(net713612), .ZN(n24349) );
  NAND2_X1 U19777 ( .A1(n24299), .A2(net742157), .ZN(n24350) );
  OR2_X1 U19778 ( .A1(n24124), .A2(n25576), .ZN(n24352) );
  CLKBUF_X1 U19779 ( .A(net713627), .Z(net749343) );
  NOR2_X1 U19780 ( .A1(n26019), .A2(n24537), .ZN(n24354) );
  NOR2_X1 U19781 ( .A1(n26019), .A2(n24537), .ZN(n24353) );
  CLKBUF_X1 U19782 ( .A(net742224), .Z(net749334) );
  OAI222_X1 U19783 ( .A1(net755757), .A2(net755238), .B1(net717055), .B2(
        net750274), .C1(net796212), .C2(net749822), .ZN(n24391) );
  INV_X1 U19784 ( .A(net750277), .ZN(net717463) );
  NOR2_X1 U19785 ( .A1(n25388), .A2(n25755), .ZN(net749312) );
  NOR3_X1 U19786 ( .A1(n25399), .A2(n25400), .A3(n25401), .ZN(net749308) );
  AND2_X1 U19787 ( .A1(n24086), .A2(net728158), .ZN(n25438) );
  CLKBUF_X1 U19788 ( .A(net714077), .Z(net749295) );
  AND2_X1 U19789 ( .A1(n24355), .A2(net713151), .ZN(n25411) );
  INV_X1 U19790 ( .A(n26055), .ZN(n25501) );
  XNOR2_X1 U19791 ( .A(n26204), .B(net716221), .ZN(n24356) );
  INV_X1 U19792 ( .A(net715048), .ZN(net749289) );
  OR2_X1 U19793 ( .A1(n25378), .A2(n25377), .ZN(n26057) );
  OR2_X1 U19794 ( .A1(n25378), .A2(n25377), .ZN(n25374) );
  INV_X1 U19795 ( .A(net736739), .ZN(net740493) );
  INV_X1 U19796 ( .A(n24358), .ZN(n24359) );
  XNOR2_X1 U19797 ( .A(n26205), .B(net716221), .ZN(n24571) );
  NOR2_X1 U19798 ( .A1(net713669), .A2(n26035), .ZN(n25938) );
  NAND2_X1 U19799 ( .A1(n25839), .A2(n25838), .ZN(n26060) );
  INV_X1 U19800 ( .A(n23993), .ZN(n25752) );
  OAI22_X1 U19801 ( .A1(n24303), .A2(net713810), .B1(net748275), .B2(net742507), .ZN(n24379) );
  INV_X1 U19802 ( .A(n26144), .ZN(n26145) );
  OR2_X1 U19803 ( .A1(n26193), .A2(n24035), .ZN(n24361) );
  INV_X1 U19804 ( .A(n26165), .ZN(n25393) );
  AND2_X1 U19805 ( .A1(DRAM_INTERFACE[0]), .A2(\core_inst/N65 ), .ZN(n297) );
  INV_X1 U19806 ( .A(net732533), .ZN(net737101) );
  AND2_X1 U19807 ( .A1(net749274), .A2(n25329), .ZN(n24376) );
  OAI22_X1 U19808 ( .A1(net737101), .A2(n4352), .B1(net741306), .B2(net738474), 
        .ZN(n25384) );
  NAND2_X1 U19809 ( .A1(net749375), .A2(n26184), .ZN(n25780) );
  INV_X1 U19810 ( .A(net717543), .ZN(net747347) );
  NOR2_X1 U19811 ( .A1(n24400), .A2(net717543), .ZN(n26172) );
  NAND2_X1 U19812 ( .A1(n24192), .A2(n24566), .ZN(n24370) );
  OAI22_X1 U19813 ( .A1(net713681), .A2(net739078), .B1(n24358), .B2(n23975), 
        .ZN(n24367) );
  OAI211_X1 U19814 ( .C1(net713677), .C2(n22673), .A(n26187), .B(n24370), .ZN(
        n24369) );
  OAI21_X1 U19815 ( .B1(net713677), .B2(net717510), .A(n24572), .ZN(n24368) );
  NAND4_X1 U19816 ( .A1(n24367), .A2(n26217), .A3(n26216), .A4(n26215), .ZN(
        n24366) );
  AOI21_X1 U19817 ( .B1(net713683), .B2(n24368), .A(n24369), .ZN(n24365) );
  NAND2_X1 U19818 ( .A1(net749832), .A2(n24170), .ZN(n24372) );
  NAND2_X1 U19819 ( .A1(n24304), .A2(n26187), .ZN(n24364) );
  AOI21_X1 U19820 ( .B1(n24365), .B2(n24366), .A(n26220), .ZN(n24363) );
  NAND4_X1 U19821 ( .A1(n24371), .A2(n24372), .A3(net713692), .A4(n24373), 
        .ZN(n24362) );
  AOI22_X1 U19822 ( .A1(n22850), .A2(n24362), .B1(n24363), .B2(n24364), .ZN(
        n26236) );
  OAI22_X1 U19823 ( .A1(net717615), .A2(net780186), .B1(net718361), .B2(n25307), .ZN(n24375) );
  NAND2_X1 U19824 ( .A1(n24356), .A2(n23969), .ZN(n25981) );
  NAND2_X1 U19825 ( .A1(net712882), .A2(n24562), .ZN(net714006) );
  NAND3_X1 U19826 ( .A1(n25382), .A2(net742286), .A3(n25423), .ZN(n25424) );
  OAI22_X1 U19827 ( .A1(n24303), .A2(net749260), .B1(n24560), .B2(net748269), 
        .ZN(n24378) );
  INV_X1 U19828 ( .A(n24378), .ZN(n25807) );
  NAND2_X1 U19829 ( .A1(net742248), .A2(net713740), .ZN(n24377) );
  OAI22_X1 U19830 ( .A1(net742508), .A2(n24303), .B1(net713851), .B2(net742259), .ZN(n25925) );
  NAND2_X1 U19831 ( .A1(net717462), .A2(net713740), .ZN(net712470) );
  MUX2_X1 U19832 ( .A(net713728), .B(net717087), .S(n24170), .Z(n24390) );
  MUX2_X1 U19833 ( .A(net713726), .B(n25662), .S(n24170), .Z(n24389) );
  MUX2_X1 U19834 ( .A(n24389), .B(n24390), .S(net750093), .Z(n24388) );
  OAI21_X1 U19835 ( .B1(net714344), .B2(net714182), .A(n24388), .ZN(n24387) );
  OAI22_X1 U19836 ( .A1(net762753), .A2(n24277), .B1(net749387), .B2(n26031), 
        .ZN(n24393) );
  OAI22_X1 U19837 ( .A1(net742483), .A2(net750287), .B1(n24560), .B2(n24358), 
        .ZN(n24392) );
  AOI22_X1 U19838 ( .A1(net767208), .A2(n24561), .B1(n26039), .B2(net714306), 
        .ZN(n24386) );
  AOI21_X1 U19839 ( .B1(net714309), .B2(n25594), .A(n24387), .ZN(n24385) );
  NOR4_X1 U19840 ( .A1(n24391), .A2(n24392), .A3(n24393), .A4(n24394), .ZN(
        n24384) );
  OAI211_X1 U19841 ( .C1(n24384), .C2(net767203), .A(n24385), .B(n24386), .ZN(
        n24383) );
  NAND2_X1 U19842 ( .A1(n24396), .A2(n24395), .ZN(n26179) );
  XNOR2_X1 U19843 ( .A(n26179), .B(net716223), .ZN(net714123) );
  NAND2_X1 U19844 ( .A1(n26180), .A2(net714123), .ZN(net714845) );
  NAND3_X1 U19845 ( .A1(n25779), .A2(net742339), .A3(n24294), .ZN(net713864)
         );
  INV_X1 U19846 ( .A(net742242), .ZN(net747343) );
  NAND2_X1 U19847 ( .A1(net747343), .A2(net715313), .ZN(n24400) );
  NAND2_X1 U19848 ( .A1(net750158), .A2(net749343), .ZN(n25773) );
  INV_X1 U19849 ( .A(n24401), .ZN(n24402) );
  OR2_X1 U19850 ( .A1(n24402), .A2(net714559), .ZN(n25404) );
  NOR3_X1 U19851 ( .A1(net749679), .A2(net748269), .A3(net714382), .ZN(n25901)
         );
  MUX2_X1 U19852 ( .A(net767234), .B(net767168), .S(n24199), .Z(n24420) );
  MUX2_X1 U19853 ( .A(net713892), .B(n26136), .S(n24199), .Z(n24421) );
  NAND3_X1 U19854 ( .A1(n24337), .A2(n25451), .A3(net713874), .ZN(n24424) );
  NAND4_X1 U19855 ( .A1(n25421), .A2(n24536), .A3(n25466), .A4(net713779), 
        .ZN(n24423) );
  OAI211_X1 U19856 ( .C1(n26135), .C2(net713897), .A(n24423), .B(n24424), .ZN(
        n24416) );
  OAI22_X1 U19857 ( .A1(net796212), .A2(net718391), .B1(net742508), .B2(n24357), .ZN(n24410) );
  NOR2_X1 U19858 ( .A1(n24410), .A2(n24411), .ZN(n24406) );
  OAI22_X1 U19859 ( .A1(n24303), .A2(net718355), .B1(net713907), .B2(net713810), .ZN(n24408) );
  NOR2_X1 U19860 ( .A1(n24408), .A2(n24409), .ZN(n24407) );
  NOR3_X1 U19861 ( .A1(n24415), .A2(n24416), .A3(n24417), .ZN(net746687) );
  OAI22_X1 U19862 ( .A1(net762754), .A2(net749454), .B1(net717055), .B2(
        net742259), .ZN(n24414) );
  INV_X1 U19863 ( .A(n24414), .ZN(n24412) );
  NAND2_X1 U19864 ( .A1(n24406), .A2(n24407), .ZN(n24405) );
  OAI21_X1 U19865 ( .B1(n24405), .B2(n24404), .A(net767221), .ZN(net746688) );
  NAND2_X1 U19866 ( .A1(net712466), .A2(net746701), .ZN(n24413) );
  NAND2_X1 U19867 ( .A1(n24418), .A2(n24419), .ZN(n24417) );
  NOR2_X1 U19868 ( .A1(net713894), .A2(net749977), .ZN(n24415) );
  OAI211_X1 U19869 ( .C1(n25599), .C2(net755699), .A(n24412), .B(n24413), .ZN(
        n24404) );
  NAND3_X1 U19870 ( .A1(n24307), .A2(n24034), .A3(net733611), .ZN(net713833)
         );
  NAND2_X1 U19871 ( .A1(net755708), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/CLA_PG_NET/N1 ), .ZN(
        n26582) );
  OAI21_X1 U19872 ( .B1(net712353), .B2(net760161), .A(n26708), .ZN(n26782) );
  NAND2_X1 U19873 ( .A1(n18398), .A2(n24731), .ZN(n24431) );
  NAND4_X1 U19874 ( .A1(n24433), .A2(n18945), .A3(n18937), .A4(n18944), .ZN(
        n24429) );
  NAND4_X1 U19875 ( .A1(n18926), .A2(n24434), .A3(n18927), .A4(n24432), .ZN(
        n24428) );
  OAI21_X1 U19876 ( .B1(n24428), .B2(n24429), .A(n25664), .ZN(n24426) );
  OAI21_X1 U19877 ( .B1(n24426), .B2(net804641), .A(n24427), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_19/N3 ) );
  NAND2_X1 U19878 ( .A1(net767238), .A2(n24732), .ZN(n24440) );
  NAND4_X1 U19879 ( .A1(n24442), .A2(n18752), .A3(n18744), .A4(n18751), .ZN(
        n24438) );
  NAND4_X1 U19880 ( .A1(n18733), .A2(n24443), .A3(n18734), .A4(n24441), .ZN(
        n24437) );
  OAI21_X1 U19881 ( .B1(n24437), .B2(n24438), .A(n26717), .ZN(n24435) );
  OAI21_X1 U19882 ( .B1(net716377), .B2(n24435), .A(n24436), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_25/N3 ) );
  NAND3_X1 U19883 ( .A1(n24460), .A2(n24461), .A3(n24462), .ZN(n24449) );
  NAND3_X1 U19884 ( .A1(n24477), .A2(n24478), .A3(n24479), .ZN(n24476) );
  NAND3_X1 U19885 ( .A1(net716261), .A2(n26670), .A3(net712397), .ZN(n24444)
         );
  NAND2_X1 U19886 ( .A1(n24445), .A2(n24444), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_28/N3 ) );
  OR2_X1 U19887 ( .A1(n24008), .A2(n24446), .ZN(n24484) );
  OR2_X1 U19888 ( .A1(net742593), .A2(n24484), .ZN(n24445) );
  NAND3_X1 U19889 ( .A1(n24488), .A2(n24489), .A3(n24490), .ZN(n24487) );
  NAND3_X1 U19890 ( .A1(n24507), .A2(n24508), .A3(n24509), .ZN(n24500) );
  NAND3_X1 U19891 ( .A1(n24513), .A2(n24514), .A3(n24515), .ZN(n24512) );
  NAND3_X1 U19892 ( .A1(n24519), .A2(n24520), .A3(n24521), .ZN(n24511) );
  NAND3_X1 U19893 ( .A1(net716261), .A2(n26327), .A3(net717049), .ZN(n24485)
         );
  NAND2_X1 U19894 ( .A1(n24485), .A2(n24486), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_16/N3 ) );
  AND2_X1 U19895 ( .A1(n25940), .A2(n25935), .ZN(n24549) );
  MUX2_X2 U19896 ( .A(n24524), .B(n25985), .S(net742092), .Z(n26135) );
  NAND2_X1 U19897 ( .A1(n24524), .A2(net742092), .ZN(n25959) );
  AND3_X1 U19898 ( .A1(n22813), .A2(n26237), .A3(n24843), .ZN(n26252) );
  INV_X1 U19899 ( .A(n26209), .ZN(n24525) );
  INV_X1 U19900 ( .A(net795568), .ZN(net716261) );
  AND2_X1 U19901 ( .A1(net742648), .A2(n24526), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_22/N3 ) );
  INV_X1 U19902 ( .A(net795568), .ZN(net742649) );
  AND2_X1 U19903 ( .A1(net716267), .A2(n18062), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_5/N3 ) );
  AND2_X1 U19904 ( .A1(net716253), .A2(n25335), .ZN(n26741) );
  INV_X1 U19905 ( .A(net765318), .ZN(net742593) );
  AND2_X1 U19906 ( .A1(net716259), .A2(n17988), .ZN(
        \core_inst/IDEX_NPC/DFF_3/N3 ) );
  AND2_X1 U19907 ( .A1(net716255), .A2(n17957), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_4/N3 ) );
  AND2_X1 U19908 ( .A1(net742648), .A2(n13778), .ZN(
        \core_inst/IDEX_NPC/DFF_12/N3 ) );
  AND2_X1 U19909 ( .A1(net742649), .A2(n17876), .ZN(
        \core_inst/IDEX_NPC/DFF_11/N3 ) );
  AND2_X1 U19910 ( .A1(net785255), .A2(n17656), .ZN(
        \core_inst/EXMEM_RF_ADDR_DEST/DFF_4/N3 ) );
  AND2_X1 U19911 ( .A1(net765318), .A2(n17654), .ZN(
        \core_inst/EXMEM_RF_ADDR_DEST/DFF_3/N3 ) );
  AND2_X1 U19912 ( .A1(net716259), .A2(n17842), .ZN(
        \core_inst/IDEX_NPC/DFF_14/N3 ) );
  AND2_X1 U19913 ( .A1(net716253), .A2(n17657), .ZN(
        \core_inst/EXMEM_RF_ADDR_DEST/DFF_2/N3 ) );
  AND2_X1 U19914 ( .A1(net716243), .A2(n17825), .ZN(
        \core_inst/IDEX_NPC/DFF_15/N3 ) );
  AND2_X1 U19915 ( .A1(net716255), .A2(n18020), .ZN(
        \core_inst/IDEX_NPC/DFF_1/N3 ) );
  AND2_X1 U19916 ( .A1(net716267), .A2(n18066), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_9/N3 ) );
  AND2_X1 U19917 ( .A1(net716259), .A2(\core_inst/s_IF_OUT_IR_OUT [0]), .ZN(
        \core_inst/IFID_IR/DFF_0/N3 ) );
  AND2_X1 U19918 ( .A1(net742649), .A2(\core_inst/s_IF_OUT_IR_OUT [10]), .ZN(
        \core_inst/IFID_IR/DFF_10/N3 ) );
  AND2_X1 U19919 ( .A1(net716267), .A2(\core_inst/s_IF_OUT_IR_OUT [13]), .ZN(
        \core_inst/IFID_IR/DFF_13/N3 ) );
  AND2_X1 U19920 ( .A1(net716267), .A2(\core_inst/s_IF_OUT_IR_OUT [16]), .ZN(
        \core_inst/IFID_IR/DFF_16/N3 ) );
  AND2_X1 U19921 ( .A1(net716267), .A2(\core_inst/s_IF_OUT_IR_OUT [1]), .ZN(
        \core_inst/IFID_IR/DFF_1/N3 ) );
  AND2_X1 U19922 ( .A1(net765341), .A2(\core_inst/s_IF_OUT_IR_OUT [3]), .ZN(
        \core_inst/IFID_IR/DFF_3/N3 ) );
  AND2_X1 U19923 ( .A1(net716267), .A2(n18056), .ZN(
        \core_inst/EXMEM_IR/DFF_14/N3 ) );
  AND2_X1 U19924 ( .A1(net741999), .A2(\core_inst/s_IF_OUT_IR_OUT [12]), .ZN(
        \core_inst/IFID_IR/DFF_12/N3 ) );
  AND2_X1 U19925 ( .A1(net716259), .A2(\core_inst/s_IF_OUT_IR_OUT [8]), .ZN(
        \core_inst/IFID_IR/DFF_8/N3 ) );
  AND2_X1 U19926 ( .A1(net765341), .A2(\core_inst/s_IF_OUT_IR_OUT [11]), .ZN(
        \core_inst/IFID_IR/DFF_11/N3 ) );
  AND2_X1 U19927 ( .A1(net742648), .A2(\core_inst/s_IF_OUT_IR_OUT [19]), .ZN(
        \core_inst/IFID_IR/DFF_19/N3 ) );
  AND2_X1 U19928 ( .A1(net742649), .A2(n18058), .ZN(
        \core_inst/EXMEM_IR/DFF_15/N3 ) );
  AND2_X1 U19929 ( .A1(net716267), .A2(n18065), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_8/N3 ) );
  AND2_X1 U19930 ( .A1(net742648), .A2(\core_inst/s_IF_OUT_IR_OUT [28]), .ZN(
        \core_inst/IFID_IR/DFF_28/N3 ) );
  AND2_X1 U19931 ( .A1(net716253), .A2(\core_inst/s_IF_OUT_IR_OUT [27]), .ZN(
        \core_inst/IFID_IR/DFF_27/N3 ) );
  AND2_X1 U19932 ( .A1(net716253), .A2(\core_inst/s_IF_OUT_IR_OUT [20]), .ZN(
        \core_inst/IFID_IR/DFF_20/N3 ) );
  AND2_X1 U19933 ( .A1(net785255), .A2(\core_inst/s_IF_OUT_IR_OUT [22]), .ZN(
        \core_inst/IFID_IR/DFF_22/N3 ) );
  AND2_X1 U19934 ( .A1(net716243), .A2(\core_inst/s_IF_OUT_IR_OUT [30]), .ZN(
        \core_inst/IFID_IR/DFF_30/N3 ) );
  INV_X1 U19935 ( .A(n26519), .ZN(\core_inst/IDEX_RF_IN1/DFF_20/N3 ) );
  INV_X1 U19936 ( .A(n26493), .ZN(\core_inst/IDEX_RF_IN2/DFF_1/N3 ) );
  INV_X1 U19937 ( .A(n26420), .ZN(\core_inst/IDEX_RF_IN1/DFF_24/N3 ) );
  INV_X1 U19938 ( .A(n26481), .ZN(\core_inst/IDEX_RF_IN1/DFF_23/N3 ) );
  INV_X1 U19939 ( .A(n26323), .ZN(\core_inst/IDEX_RF_IN2/DFF_0/N3 ) );
  INV_X1 U19940 ( .A(n26713), .ZN(n11847) );
  INV_X1 U19941 ( .A(n25852), .ZN(n25442) );
  OR2_X1 U19942 ( .A1(net713602), .A2(n25944), .ZN(n24528) );
  NOR2_X1 U19943 ( .A1(n24319), .A2(n24089), .ZN(n24529) );
  BUF_X2 U19944 ( .A(net713560), .Z(net742508) );
  OR2_X1 U19945 ( .A1(n25405), .A2(n25874), .ZN(n24530) );
  INV_X1 U19946 ( .A(net713607), .ZN(net713560) );
  OR2_X1 U19947 ( .A1(net718134), .A2(n24786), .ZN(n25385) );
  AND2_X1 U19948 ( .A1(net740526), .A2(net755714), .ZN(net734385) );
  CLKBUF_X1 U19949 ( .A(net713677), .Z(net742483) );
  INV_X1 U19950 ( .A(net713905), .ZN(net742473) );
  CLKBUF_X1 U19951 ( .A(n26089), .Z(n24532) );
  INV_X1 U19952 ( .A(n24531), .ZN(n25816) );
  INV_X1 U19953 ( .A(n24307), .ZN(n25437) );
  AOI22_X1 U19954 ( .A1(n26137), .A2(net713779), .B1(net713870), .B2(net713874), .ZN(n24533) );
  CLKBUF_X1 U19955 ( .A(n26726), .Z(n24534) );
  NOR2_X1 U19956 ( .A1(n25805), .A2(n25804), .ZN(n26726) );
  INV_X1 U19957 ( .A(n24282), .ZN(n25874) );
  INV_X1 U19958 ( .A(net734607), .ZN(net712378) );
  CLKBUF_X1 U19959 ( .A(net715443), .Z(net742412) );
  INV_X1 U19960 ( .A(net750135), .ZN(net742413) );
  INV_X1 U19961 ( .A(n26711), .ZN(n14058) );
  INV_X1 U19962 ( .A(n26716), .ZN(n11725) );
  INV_X1 U19963 ( .A(net718103), .ZN(net714611) );
  INV_X1 U19964 ( .A(net712879), .ZN(net713167) );
  INV_X1 U19965 ( .A(net712384), .ZN(net712344) );
  AND2_X1 U19966 ( .A1(net716259), .A2(s_IFID_IR[30]), .ZN(
        \core_inst/IDEX_IR/DFF_30/N3 ) );
  INV_X1 U19967 ( .A(n26708), .ZN(\core_inst/IFID_NPC/DFF_12/N3 ) );
  INV_X1 U19968 ( .A(n26712), .ZN(\core_inst/IFID_NPC/DFF_16/N3 ) );
  INV_X1 U19969 ( .A(n26719), .ZN(n15062) );
  OR2_X1 U19970 ( .A1(n25454), .A2(n25456), .ZN(n25315) );
  INV_X1 U19971 ( .A(net714551), .ZN(net740526) );
  AND2_X1 U19972 ( .A1(n24296), .A2(net750019), .ZN(n24537) );
  INV_X1 U19973 ( .A(net713707), .ZN(net742325) );
  INV_X1 U19974 ( .A(net713707), .ZN(net742324) );
  INV_X1 U19975 ( .A(net713707), .ZN(net713701) );
  INV_X1 U19976 ( .A(n24333), .ZN(n24538) );
  OAI21_X1 U19977 ( .B1(n25855), .B2(n26072), .A(n25976), .ZN(net742309) );
  OAI21_X1 U19978 ( .B1(n25855), .B2(n26072), .A(n25976), .ZN(n26119) );
  INV_X1 U19979 ( .A(net714977), .ZN(net714855) );
  INV_X1 U19980 ( .A(n26071), .ZN(n24539) );
  INV_X1 U19981 ( .A(net749707), .ZN(net714007) );
  CLKBUF_X1 U19982 ( .A(net714076), .Z(net742296) );
  CLKBUF_X1 U19983 ( .A(n26088), .Z(n24540) );
  INV_X1 U19984 ( .A(net749725), .ZN(net713679) );
  MUX2_X2 U19985 ( .A(n869), .B(n26089), .S(net787526), .Z(net713612) );
  INV_X1 U19986 ( .A(net717103), .ZN(net713845) );
  AND2_X2 U19987 ( .A1(n24268), .A2(n24608), .ZN(n24543) );
  OR2_X1 U19988 ( .A1(net716237), .A2(\core_inst/EXMEM_NPC/DFF_18/N3 ), .ZN(
        n24608) );
  NOR2_X1 U19989 ( .A1(net742243), .A2(net749273), .ZN(net742248) );
  NOR2_X1 U19990 ( .A1(net796014), .A2(net742243), .ZN(n25417) );
  INV_X1 U19991 ( .A(n26140), .ZN(n26142) );
  INV_X1 U19992 ( .A(n26022), .ZN(n26027) );
  INV_X1 U19993 ( .A(n26561), .ZN(n25365) );
  BUF_X2 U19994 ( .A(n25443), .Z(n24546) );
  NAND2_X1 U19995 ( .A1(net749372), .A2(net713733), .ZN(n25443) );
  INV_X1 U19996 ( .A(net714401), .ZN(net713979) );
  OR2_X1 U19997 ( .A1(n25782), .A2(net717511), .ZN(n25600) );
  INV_X1 U19998 ( .A(n25782), .ZN(n25786) );
  NAND3_X1 U19999 ( .A1(n24314), .A2(n25510), .A3(n25511), .ZN(n24551) );
  INV_X1 U20000 ( .A(n25972), .ZN(n25973) );
  OR3_X1 U20001 ( .A1(n25441), .A2(n25439), .A3(n25440), .ZN(n24553) );
  INV_X1 U20002 ( .A(net713687), .ZN(net713754) );
  AND2_X1 U20003 ( .A1(n26151), .A2(n25579), .ZN(n26152) );
  NOR2_X1 U20004 ( .A1(net767203), .A2(n24175), .ZN(n25989) );
  NOR2_X1 U20005 ( .A1(n25393), .A2(n24298), .ZN(net713740) );
  INV_X1 U20006 ( .A(n26149), .ZN(n24555) );
  INV_X1 U20007 ( .A(n26149), .ZN(n24554) );
  CLKBUF_X1 U20008 ( .A(n26061), .Z(n24556) );
  INV_X1 U20009 ( .A(net713811), .ZN(net713964) );
  BUF_X1 U20010 ( .A(n25418), .Z(n24558) );
  NOR2_X1 U20011 ( .A1(n25577), .A2(n24271), .ZN(net715284) );
  OR2_X1 U20012 ( .A1(net715359), .A2(n24266), .ZN(n24559) );
  INV_X1 U20013 ( .A(net713740), .ZN(net715359) );
  INV_X1 U20014 ( .A(n26063), .ZN(n25412) );
  INV_X1 U20015 ( .A(net713733), .ZN(net737907) );
  INV_X1 U20016 ( .A(net714602), .ZN(net714585) );
  INV_X1 U20017 ( .A(net749372), .ZN(net713990) );
  INV_X1 U20018 ( .A(n25443), .ZN(n25467) );
  NOR2_X1 U20019 ( .A1(net750019), .A2(n24296), .ZN(n26118) );
  INV_X1 U20020 ( .A(net713985), .ZN(net713867) );
  XNOR2_X1 U20021 ( .A(n25579), .B(net716215), .ZN(n24564) );
  INV_X1 U20022 ( .A(net755258), .ZN(net714871) );
  INV_X1 U20023 ( .A(net749830), .ZN(net742061) );
  INV_X1 U20024 ( .A(n26077), .ZN(n26079) );
  INV_X1 U20025 ( .A(net742265), .ZN(net715422) );
  INV_X1 U20026 ( .A(net742046), .ZN(net742047) );
  INV_X1 U20027 ( .A(net712882), .ZN(net715048) );
  INV_X1 U20028 ( .A(n26105), .ZN(n26109) );
  INV_X1 U20029 ( .A(n25835), .ZN(n25514) );
  INV_X1 U20030 ( .A(net750277), .ZN(net717462) );
  NAND2_X1 U20031 ( .A1(net749307), .A2(net786867), .ZN(n24568) );
  AND2_X1 U20032 ( .A1(net742368), .A2(n17792), .ZN(
        \core_inst/IDEX_NPC/DFF_16/N3 ) );
  AND2_X1 U20033 ( .A1(net716265), .A2(n17736), .ZN(
        \core_inst/IDEX_NPC/DFF_24/N3 ) );
  AND2_X1 U20034 ( .A1(net716385), .A2(n17707), .ZN(
        \core_inst/IDEX_NPC/DFF_30/N3 ) );
  AND2_X1 U20035 ( .A1(net716257), .A2(n17778), .ZN(
        \core_inst/IDEX_NPC/DFF_19/N3 ) );
  AND2_X1 U20036 ( .A1(net716243), .A2(n17764), .ZN(
        \core_inst/IDEX_NPC/DFF_22/N3 ) );
  AND2_X1 U20037 ( .A1(net742649), .A2(n17700), .ZN(
        \core_inst/IDEX_NPC/DFF_31/N3 ) );
  AND2_X1 U20038 ( .A1(net716255), .A2(n18054), .ZN(
        \core_inst/EXMEM_IR/DFF_11/N3 ) );
  AND2_X1 U20039 ( .A1(net742648), .A2(n17696), .ZN(
        \core_inst/IDEX_NPC/DFF_29/N3 ) );
  AND2_X1 U20040 ( .A1(net742649), .A2(n17744), .ZN(
        \core_inst/IDEX_NPC/DFF_17/N3 ) );
  AND2_X1 U20041 ( .A1(net716253), .A2(n18063), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_6/N3 ) );
  AND2_X1 U20042 ( .A1(net742648), .A2(n18064), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_7/N3 ) );
  AND2_X1 U20043 ( .A1(net716255), .A2(n17808), .ZN(
        \core_inst/IDEX_NPC/DFF_13/N3 ) );
  AND2_X1 U20044 ( .A1(net742649), .A2(n17771), .ZN(
        \core_inst/IDEX_NPC/DFF_20/N3 ) );
  AND2_X1 U20045 ( .A1(net716385), .A2(n17729), .ZN(
        \core_inst/IDEX_NPC/DFF_26/N3 ) );
  OR2_X1 U20046 ( .A1(net765629), .A2(n22677), .ZN(net724631) );
  INV_X1 U20047 ( .A(n25751), .ZN(n25748) );
  OR2_X1 U20048 ( .A1(net767341), .A2(n6156), .ZN(net724630) );
  NOR2_X1 U20049 ( .A1(n24276), .A2(net796258), .ZN(n24570) );
  AND2_X1 U20050 ( .A1(net716243), .A2(\core_inst/s_IF_OUT_IR_OUT [18]), .ZN(
        \core_inst/IFID_IR/DFF_18/N3 ) );
  INV_X1 U20051 ( .A(net717059), .ZN(net712467) );
  INV_X1 U20052 ( .A(n24552), .ZN(n25999) );
  INV_X1 U20053 ( .A(net742284), .ZN(net715421) );
  AND2_X1 U20054 ( .A1(n25423), .A2(n25382), .ZN(n26034) );
  INV_X1 U20055 ( .A(net749292), .ZN(net712356) );
  INV_X1 U20056 ( .A(n26019), .ZN(n25971) );
  INV_X1 U20057 ( .A(n26212), .ZN(n25909) );
  INV_X1 U20058 ( .A(net749566), .ZN(net712390) );
  INV_X1 U20059 ( .A(net715614), .ZN(net715615) );
  CLKBUF_X3 U20060 ( .A(n26065), .Z(n24577) );
  INV_X1 U20061 ( .A(n26042), .ZN(n26065) );
  INV_X1 U20062 ( .A(n24566), .ZN(n25413) );
  AND2_X1 U20063 ( .A1(net713454), .A2(n24291), .ZN(n26120) );
  INV_X1 U20064 ( .A(n23027), .ZN(n26114) );
  INV_X1 U20065 ( .A(n25390), .ZN(n25391) );
  INV_X1 U20066 ( .A(n26180), .ZN(n26071) );
  NOR2_X1 U20067 ( .A1(n26058), .A2(n24312), .ZN(n26214) );
  INV_X1 U20068 ( .A(net713677), .ZN(net714194) );
  NAND2_X1 U20069 ( .A1(net713677), .A2(n24281), .ZN(net714977) );
  INV_X1 U20070 ( .A(n25418), .ZN(n25815) );
  AND2_X1 U20071 ( .A1(net749507), .A2(net749428), .ZN(n25598) );
  INV_X1 U20072 ( .A(n26404), .ZN(n25597) );
  AND2_X1 U20073 ( .A1(n24098), .A2(net734022), .ZN(n25406) );
  INV_X1 U20074 ( .A(n24570), .ZN(n25599) );
  INV_X1 U20075 ( .A(net742309), .ZN(net712872) );
  MUX2_X2 U20076 ( .A(\core_inst/EXMEM_NPC/DFF_29/N3 ), .B(n26107), .S(
        net716237), .Z(net713985) );
  INV_X1 U20077 ( .A(net713627), .ZN(net713633) );
  OR2_X1 U20078 ( .A1(net749525), .A2(n24531), .ZN(n24843) );
  AND2_X1 U20079 ( .A1(net749525), .A2(n26143), .ZN(n26146) );
  AND3_X1 U20080 ( .A1(n24283), .A2(net742326), .A3(net733611), .ZN(n26404) );
  INV_X1 U20081 ( .A(net713570), .ZN(net731327) );
  MUX2_X2 U20082 ( .A(\core_inst/EXMEM_NPC/DFF_10/N3 ), .B(n26111), .S(
        net716237), .Z(net713707) );
  INV_X1 U20083 ( .A(n24565), .ZN(n25994) );
  INV_X1 U20084 ( .A(n24338), .ZN(n25402) );
  INV_X2 U20085 ( .A(net749993), .ZN(net713753) );
  INV_X1 U20086 ( .A(net717053), .ZN(net712466) );
  BUF_X2 U20087 ( .A(net717720), .Z(net718341) );
  INV_X1 U20088 ( .A(net715632), .ZN(net715460) );
  INV_X1 U20089 ( .A(net750228), .ZN(net713711) );
  OR2_X1 U20090 ( .A1(n25398), .A2(n26070), .ZN(n25423) );
  AND2_X1 U20091 ( .A1(net716243), .A2(\core_inst/s_IF_OUT_IR_OUT [9]), .ZN(
        \core_inst/IFID_IR/DFF_9/N3 ) );
  AND2_X1 U20092 ( .A1(net785255), .A2(\core_inst/s_IF_OUT_IR_OUT [7]), .ZN(
        \core_inst/IFID_IR/DFF_7/N3 ) );
  AND2_X1 U20093 ( .A1(net716263), .A2(\core_inst/s_IF_OUT_IR_OUT [5]), .ZN(
        \core_inst/IFID_IR/DFF_5/N3 ) );
  AND2_X1 U20094 ( .A1(net742576), .A2(\core_inst/s_IF_OUT_IR_OUT [25]), .ZN(
        \core_inst/IFID_IR/DFF_25/N3 ) );
  AND2_X1 U20095 ( .A1(net716253), .A2(\core_inst/s_IF_OUT_IR_OUT [4]), .ZN(
        \core_inst/IFID_IR/DFF_4/N3 ) );
  NAND2_X1 U20096 ( .A1(n24299), .A2(net742157), .ZN(n25940) );
  INV_X1 U20097 ( .A(n26149), .ZN(n26058) );
  AND2_X1 U20098 ( .A1(net716265), .A2(\core_inst/s_IF_OUT_IR_OUT [15]), .ZN(
        \core_inst/IFID_IR/DFF_15/N3 ) );
  AND2_X1 U20099 ( .A1(net765341), .A2(\core_inst/s_IF_OUT_IR_OUT [6]), .ZN(
        \core_inst/IFID_IR/DFF_6/N3 ) );
  AND2_X1 U20100 ( .A1(net742576), .A2(\core_inst/s_IF_OUT_IR_OUT [24]), .ZN(
        \core_inst/IFID_IR/DFF_24/N3 ) );
  AND2_X1 U20101 ( .A1(net741999), .A2(\core_inst/s_IF_OUT_IR_OUT [31]), .ZN(
        \core_inst/IFID_IR/DFF_31/N3 ) );
  AND2_X1 U20102 ( .A1(net716385), .A2(\core_inst/s_IF_OUT_IR_OUT [17]), .ZN(
        \core_inst/IFID_IR/DFF_17/N3 ) );
  INV_X1 U20103 ( .A(net750135), .ZN(net715419) );
  INV_X1 U20104 ( .A(net750135), .ZN(net718432) );
  INV_X1 U20105 ( .A(net750135), .ZN(net718154) );
  NOR2_X1 U20106 ( .A1(net796193), .A2(n6562), .ZN(n26743) );
  NOR2_X1 U20107 ( .A1(net796193), .A2(n5611), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_12/N3 ) );
  NOR2_X1 U20108 ( .A1(net796143), .A2(n22675), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_20/N3 ) );
  NOR2_X1 U20109 ( .A1(net796143), .A2(n22676), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_18/N3 ) );
  NOR2_X1 U20110 ( .A1(net812279), .A2(n1301), .ZN(
        \core_inst/IDEX_NPC/DFF_7/N3 ) );
  NOR2_X1 U20111 ( .A1(net716367), .A2(net780188), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_3/N3 ) );
  NOR2_X1 U20112 ( .A1(net796193), .A2(n25322), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_8/N3 ) );
  NOR2_X1 U20113 ( .A1(net796137), .A2(n24610), .ZN(n26781) );
  NOR2_X1 U20114 ( .A1(net796136), .A2(net717952), .ZN(
        \core_inst/EXMEM_IR/DFF_18/N3 ) );
  AOI21_X1 U20115 ( .B1(n26626), .B2(n26625), .A(net716331), .ZN(
        \core_inst/IDEX_RF_IN1/DFF_3/N3 ) );
  AOI21_X1 U20116 ( .B1(n25524), .B2(n25525), .A(net796232), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_2/N3 ) );
  AOI21_X1 U20117 ( .B1(n25516), .B2(n25517), .A(net796143), .ZN(
        \core_inst/IDEX_RF_IN1/DFF_4/N3 ) );
  AOI21_X1 U20118 ( .B1(n25532), .B2(n25533), .A(net796232), .ZN(
        \core_inst/IDEX_RF_IN1/DFF_8/N3 ) );
  NOR2_X1 U20119 ( .A1(net716367), .A2(n1668), .ZN(
        \core_inst/EXMEM_IR/DFF_19/N3 ) );
  NOR2_X1 U20120 ( .A1(net716311), .A2(n24585), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_3/N3 ) );
  AOI21_X1 U20121 ( .B1(n26545), .B2(n26544), .A(net796232), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_7/N3 ) );
  AOI21_X1 U20122 ( .B1(n26373), .B2(n26372), .A(net716369), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_3/N3 ) );
  AOI21_X1 U20123 ( .B1(n26290), .B2(n26289), .A(net796232), .ZN(
        \core_inst/IDEX_RF_IN1/DFF_13/N3 ) );
  AOI21_X1 U20124 ( .B1(n26621), .B2(n26620), .A(net716377), .ZN(
        \core_inst/IDEX_RF_IN1/DFF_2/N3 ) );
  AOI21_X1 U20125 ( .B1(n26557), .B2(n26556), .A(net716333), .ZN(
        \core_inst/IDEX_RF_IN1/DFF_5/N3 ) );
  AOI21_X1 U20126 ( .B1(n26504), .B2(n26503), .A(net796136), .ZN(
        \core_inst/IDEX_RF_IN1/DFF_6/N3 ) );
  AOI21_X1 U20127 ( .B1(n26344), .B2(n26343), .A(net796143), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_8/N3 ) );
  NOR2_X1 U20128 ( .A1(net812279), .A2(net741576), .ZN(
        \core_inst/EXMEM_IR/DFF_26/N3 ) );
  NAND2_X1 U20129 ( .A1(n26457), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [26]), .ZN(n26558) );
  NAND2_X1 U20130 ( .A1(n26570), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [24]), .ZN(net712838) );
  NAND2_X1 U20131 ( .A1(n26579), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [16]), .ZN(n26578) );
  NAND2_X1 U20132 ( .A1(net712488), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [14]), .ZN(net712490) );
  NAND2_X1 U20133 ( .A1(n26575), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [10]), .ZN(n26459) );
  NAND2_X1 U20134 ( .A1(n26572), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [8]), .ZN(n26576) );
  NAND2_X1 U20135 ( .A1(n26709), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [6]), .ZN(n26671) );
  NAND2_X1 U20136 ( .A1(n26604), .A2(
        \core_inst/IF_stage/PLUS4_ADDER/CARRY_GENERATOR/s_CLA_CGEN_pg_network_p [4]), .ZN(n26710) );
  NAND2_X1 U20137 ( .A1(n24542), .A2(n26246), .ZN(n26249) );
  NAND2_X1 U20138 ( .A1(n26231), .A2(n26232), .ZN(n26241) );
  NAND2_X1 U20139 ( .A1(net749454), .A2(n26208), .ZN(n26207) );
  NAND2_X1 U20140 ( .A1(n26038), .A2(net749732), .ZN(n25410) );
  NAND4_X1 U20141 ( .A1(n26176), .A2(n26177), .A3(n23975), .A4(n26178), .ZN(
        n25409) );
  NAND2_X1 U20142 ( .A1(n26173), .A2(net750264), .ZN(n26177) );
  NOR2_X1 U20143 ( .A1(n26240), .A2(net713728), .ZN(net713763) );
  AOI21_X1 U20144 ( .B1(n26167), .B2(n26166), .A(n25380), .ZN(net713761) );
  AOI21_X1 U20145 ( .B1(n26163), .B2(net713779), .A(n26162), .ZN(n26167) );
  NOR3_X1 U20146 ( .A1(n26161), .A2(n26160), .A3(n26159), .ZN(n26162) );
  NAND2_X1 U20147 ( .A1(n26156), .A2(n26155), .ZN(n26160) );
  NOR2_X1 U20148 ( .A1(n25471), .A2(n25467), .ZN(net713857) );
  NOR2_X1 U20149 ( .A1(n25597), .A2(net713167), .ZN(net713952) );
  NOR2_X1 U20150 ( .A1(n25598), .A2(n24191), .ZN(n26073) );
  NAND2_X1 U20151 ( .A1(net713867), .A2(n26052), .ZN(n26227) );
  NAND2_X1 U20152 ( .A1(n26071), .A2(n24171), .ZN(net713692) );
  NOR2_X1 U20153 ( .A1(n26033), .A2(n26032), .ZN(net714347) );
  NOR2_X1 U20154 ( .A1(n26030), .A2(n26029), .ZN(net714346) );
  NAND2_X1 U20155 ( .A1(net732754), .A2(net767221), .ZN(net729186) );
  NAND2_X1 U20156 ( .A1(net714559), .A2(n25990), .ZN(n26229) );
  NOR4_X1 U20157 ( .A1(n24562), .A2(n25984), .A3(net760144), .A4(net749707), 
        .ZN(n25975) );
  NAND2_X1 U20158 ( .A1(n24172), .A2(n25973), .ZN(n25984) );
  NAND2_X1 U20159 ( .A1(n26012), .A2(net366451), .ZN(net714465) );
  NOR2_X1 U20160 ( .A1(n26009), .A2(net714476), .ZN(net714464) );
  INV_X2 U20161 ( .A(net713897), .ZN(net713785) );
  BUF_X1 U20162 ( .A(net712879), .Z(net718400) );
  NOR4_X1 U20163 ( .A1(n25951), .A2(n25950), .A3(n25949), .A4(n25948), .ZN(
        n25956) );
  XNOR2_X1 U20164 ( .A(n25945), .B(net755740), .ZN(net714105) );
  NAND3_X1 U20165 ( .A1(n26074), .A2(net714104), .A3(n24191), .ZN(n26075) );
  NAND2_X1 U20166 ( .A1(net749476), .A2(net714113), .ZN(n26074) );
  OAI21_X1 U20167 ( .B1(n25897), .B2(net713154), .A(n25896), .ZN(net712445) );
  NOR4_X1 U20168 ( .A1(n25895), .A2(n25894), .A3(n25893), .A4(n25892), .ZN(
        n25896) );
  NOR2_X1 U20169 ( .A1(n26057), .A2(net714182), .ZN(n25892) );
  OAI211_X1 U20170 ( .C1(net714354), .C2(net714267), .A(n25891), .B(n25890), 
        .ZN(n25894) );
  XNOR2_X1 U20171 ( .A(n25983), .B(n25876), .ZN(n25897) );
  NAND2_X1 U20172 ( .A1(n25939), .A2(net714907), .ZN(n25983) );
  NOR2_X1 U20173 ( .A1(n25919), .A2(n25918), .ZN(net712493) );
  NOR2_X1 U20174 ( .A1(n25885), .A2(n25886), .ZN(n26028) );
  OAI21_X1 U20175 ( .B1(n24346), .B2(n26041), .A(n24197), .ZN(n26068) );
  NOR2_X1 U20176 ( .A1(n25427), .A2(net714770), .ZN(net738840) );
  AOI21_X1 U20177 ( .B1(net742146), .B2(net755139), .A(n25938), .ZN(net728823)
         );
  NAND2_X1 U20178 ( .A1(n26562), .A2(net713751), .ZN(n25875) );
  NOR2_X1 U20179 ( .A1(n26130), .A2(n26128), .ZN(n26562) );
  NAND2_X1 U20180 ( .A1(n26565), .A2(n26127), .ZN(n26130) );
  NAND2_X1 U20181 ( .A1(n25872), .A2(net713868), .ZN(n26565) );
  NAND2_X1 U20182 ( .A1(net713985), .A2(n24179), .ZN(n25873) );
  NAND2_X1 U20183 ( .A1(net767206), .A2(n25871), .ZN(n26127) );
  NAND2_X1 U20184 ( .A1(net712467), .A2(net713775), .ZN(n26055) );
  NAND3_X1 U20185 ( .A1(net726959), .A2(n25472), .A3(net726961), .ZN(n25373)
         );
  NAND2_X1 U20186 ( .A1(n25848), .A2(n25847), .ZN(n26198) );
  NAND2_X1 U20187 ( .A1(n25852), .A2(net713636), .ZN(n26021) );
  XNOR2_X1 U20188 ( .A(n26197), .B(net716223), .ZN(n25852) );
  NAND2_X1 U20189 ( .A1(n24035), .A2(n24301), .ZN(n26041) );
  NOR2_X1 U20190 ( .A1(n25842), .A2(n25841), .ZN(n25843) );
  XNOR2_X1 U20191 ( .A(n26060), .B(net716215), .ZN(n25840) );
  NAND2_X1 U20192 ( .A1(net714544), .A2(n25992), .ZN(n25515) );
  AOI21_X1 U20193 ( .B1(net713966), .B2(net714934), .A(n23023), .ZN(n25405) );
  NAND2_X1 U20194 ( .A1(n25514), .A2(n25578), .ZN(n25993) );
  NAND3_X1 U20195 ( .A1(net724630), .A2(net724632), .A3(net724631), .ZN(
        net713934) );
  NAND2_X1 U20196 ( .A1(n26564), .A2(n26119), .ZN(net714934) );
  NAND2_X1 U20197 ( .A1(n22845), .A2(net713602), .ZN(n25976) );
  NOR2_X1 U20198 ( .A1(n25944), .A2(net713602), .ZN(n25855) );
  XNOR2_X1 U20199 ( .A(n25832), .B(net716215), .ZN(n25944) );
  NOR2_X1 U20200 ( .A1(net714559), .A2(n25833), .ZN(n25834) );
  XNOR2_X1 U20201 ( .A(n25991), .B(net716215), .ZN(n25833) );
  XNOR2_X1 U20202 ( .A(n26181), .B(net716223), .ZN(net714440) );
  NAND2_X1 U20203 ( .A1(n23978), .A2(net749410), .ZN(net714287) );
  NOR2_X1 U20204 ( .A1(net750274), .A2(net755210), .ZN(n25898) );
  NOR2_X1 U20205 ( .A1(n26064), .A2(n25816), .ZN(n26186) );
  NOR2_X1 U20206 ( .A1(net715236), .A2(net715235), .ZN(n25594) );
  NOR2_X1 U20207 ( .A1(n25793), .A2(net749725), .ZN(n25513) );
  NAND3_X1 U20208 ( .A1(n24314), .A2(n25510), .A3(n25511), .ZN(n25795) );
  BUF_X1 U20209 ( .A(net713612), .Z(net718380) );
  NAND2_X1 U20210 ( .A1(n25452), .A2(n25453), .ZN(n25512) );
  NAND2_X1 U20211 ( .A1(n25449), .A2(net732762), .ZN(n25453) );
  NOR2_X1 U20212 ( .A1(n25922), .A2(n25412), .ZN(net713454) );
  NOR2_X1 U20213 ( .A1(net750024), .A2(n26061), .ZN(n26532) );
  NOR2_X1 U20214 ( .A1(n25455), .A2(n25315), .ZN(n25452) );
  NOR3_X1 U20215 ( .A1(n25441), .A2(n25439), .A3(n25440), .ZN(n26090) );
  NAND2_X1 U20216 ( .A1(n25989), .A2(net718367), .ZN(net714382) );
  OAI22_X1 U20217 ( .A1(net718154), .A2(n1740), .B1(net718337), .B2(n25312), 
        .ZN(n25763) );
  NAND2_X1 U20218 ( .A1(n26113), .A2(net716237), .ZN(n25367) );
  NOR3_X1 U20219 ( .A1(n25401), .A2(n25399), .A3(n25400), .ZN(n26078) );
  NOR2_X1 U20220 ( .A1(net715551), .A2(n25469), .ZN(n26110) );
  OAI22_X1 U20221 ( .A1(n4410), .A2(net718337), .B1(net742413), .B2(n1744), 
        .ZN(n25469) );
  NAND2_X1 U20222 ( .A1(n25989), .A2(net739078), .ZN(net713882) );
  NAND2_X1 U20223 ( .A1(net713777), .A2(n25832), .ZN(n26211) );
  OAI21_X1 U20224 ( .B1(n25457), .B2(net713751), .A(n25458), .ZN(n25455) );
  NOR4_X1 U20225 ( .A1(n25462), .A2(n25464), .A3(n25463), .A4(n25465), .ZN(
        n25457) );
  NOR2_X1 U20226 ( .A1(n25393), .A2(n24271), .ZN(net715313) );
  AND2_X2 U20227 ( .A1(n24271), .A2(n25393), .ZN(net713733) );
  OAI22_X1 U20228 ( .A1(n25595), .A2(n4421), .B1(n1750), .B2(net765744), .ZN(
        n25755) );
  NAND2_X1 U20229 ( .A1(net713845), .A2(\core_inst/MEMWB_ALUOUT/DFF_4/N3 ), 
        .ZN(n25760) );
  NAND2_X1 U20230 ( .A1(n23993), .A2(net366126), .ZN(n25507) );
  NAND3_X1 U20231 ( .A1(n25592), .A2(n25589), .A3(net718006), .ZN(n25370) );
  NAND2_X1 U20232 ( .A1(net718070), .A2(net718069), .ZN(n25746) );
  NAND2_X1 U20233 ( .A1(n25581), .A2(net334510), .ZN(n25747) );
  OAI211_X1 U20234 ( .C1(net742047), .C2(net749987), .A(net715795), .B(
        net715796), .ZN(n25751) );
  NAND3_X1 U20235 ( .A1(net715794), .A2(n24316), .A3(net742047), .ZN(net715796) );
  NOR2_X1 U20236 ( .A1(net742157), .A2(n26060), .ZN(n26190) );
  NOR2_X1 U20237 ( .A1(n24356), .A2(n23969), .ZN(n25941) );
  NAND2_X1 U20238 ( .A1(n24349), .A2(n25980), .ZN(n25942) );
  NOR2_X1 U20239 ( .A1(s_IFID_IR[21]), .A2(s_IFID_IR[25]), .ZN(n20061) );
  NAND2_X1 U20240 ( .A1(s_IFID_IR[21]), .A2(s_IFID_IR[25]), .ZN(n20068) );
  NAND2_X1 U20241 ( .A1(net715584), .A2(net741282), .ZN(n25662) );
  NOR2_X1 U20242 ( .A1(n25391), .A2(n25356), .ZN(n25439) );
  NAND2_X1 U20243 ( .A1(net715584), .A2(net741603), .ZN(net713770) );
  NOR2_X1 U20244 ( .A1(n20200), .A2(n20201), .ZN(n20183) );
  NOR2_X1 U20245 ( .A1(n20154), .A2(n20182), .ZN(n20155) );
  NOR2_X1 U20246 ( .A1(n20153), .A2(n20154), .ZN(n20134) );
  NOR2_X1 U20247 ( .A1(n20240), .A2(n20431), .ZN(n20443) );
  NOR2_X1 U20248 ( .A1(n20332), .A2(n20431), .ZN(n20501) );
  NOR2_X1 U20249 ( .A1(n20372), .A2(n20431), .ZN(n20519) );
  NOR2_X1 U20250 ( .A1(n20182), .A2(n20431), .ZN(n20581) );
  NOR2_X1 U20251 ( .A1(n20153), .A2(n20431), .ZN(n20547) );
  NOR2_X1 U20252 ( .A1(n20332), .A2(n20293), .ZN(n20367) );
  NOR2_X1 U20253 ( .A1(n20240), .A2(n20293), .ZN(n20333) );
  NOR2_X1 U20254 ( .A1(n20260), .A2(n20293), .ZN(n20350) );
  NOR2_X1 U20255 ( .A1(n20153), .A2(n20293), .ZN(n20373) );
  NOR2_X1 U20256 ( .A1(n20182), .A2(n20293), .ZN(n20392) );
  NOR2_X1 U20257 ( .A1(n20154), .A2(n20372), .ZN(n20684) );
  INV_X2 U20258 ( .A(n298), .ZN(n25684) );
  BUF_X1 U20259 ( .A(n19335), .Z(n25681) );
  BUF_X1 U20260 ( .A(n18328), .Z(net716423) );
  NOR2_X2 U20261 ( .A1(net708964), .A2(n19243), .ZN(n18373) );
  NOR2_X2 U20262 ( .A1(n19243), .A2(n19246), .ZN(n18372) );
  INV_X2 U20263 ( .A(n24615), .ZN(n25683) );
  BUF_X1 U20264 ( .A(n19393), .Z(n25674) );
  BUF_X1 U20265 ( .A(n19333), .Z(n25682) );
  NOR2_X2 U20266 ( .A1(n20069), .A2(n20067), .ZN(n19333) );
  INV_X2 U20267 ( .A(n24617), .ZN(n25678) );
  INV_X2 U20268 ( .A(n24619), .ZN(n25677) );
  NOR2_X2 U20269 ( .A1(n20081), .A2(n20069), .ZN(n19348) );
  NOR2_X2 U20270 ( .A1(n26778), .A2(n20065), .ZN(n19373) );
  NOR2_X2 U20271 ( .A1(n20065), .A2(n20068), .ZN(n19372) );
  INV_X2 U20272 ( .A(n19366), .ZN(n19336) );
  NAND2_X2 U20273 ( .A1(n25744), .A2(n20076), .ZN(n26785) );
  MUX2_X2 U20274 ( .A(n1456), .B(n26100), .S(net787512), .Z(net713677) );
  AOI22_X1 U20275 ( .A1(n20134), .A2(n26715), .B1(n25672), .B2(n3004), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_9/DFF_12/N3 ) );
  AOI22_X1 U20276 ( .A1(n20155), .A2(n26715), .B1(n25670), .B2(n24822), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_8/DFF_12/N3 ) );
  AOI22_X1 U20277 ( .A1(n20183), .A2(n26715), .B1(n25668), .B2(n24829), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_7/DFF_12/N3 ) );
  AOI22_X1 U20278 ( .A1(n24009), .A2(n26715), .B1(n20371), .B2(n24621), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_26/DFF_12/N3 ) );
  AOI22_X1 U20279 ( .A1(n24025), .A2(n26715), .B1(n20263), .B2(n24828), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_31/DFF_12/N3 ) );
  AOI22_X1 U20280 ( .A1(n24006), .A2(n26715), .B1(n20334), .B2(n24821), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_29/DFF_12/N3 ) );
  AOI22_X1 U20281 ( .A1(n24000), .A2(n26715), .B1(n20521), .B2(n24824), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_18/DFF_12/N3 ) );
  AOI22_X1 U20282 ( .A1(n23998), .A2(n26715), .B1(n20582), .B2(n24842), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_16/DFF_12/N3 ) );
  AOI22_X1 U20283 ( .A1(n24012), .A2(n26715), .B1(n20593), .B2(n24823), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_15/DFF_12/N3 ) );
  AOI22_X1 U20284 ( .A1(n24010), .A2(n26715), .B1(n20400), .B2(n24826), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_23/DFF_12/N3 ) );
  AOI22_X1 U20285 ( .A1(n24013), .A2(n26715), .B1(n20651), .B2(n24831), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_12/DFF_12/N3 ) );
  AOI22_X1 U20286 ( .A1(n24023), .A2(n26715), .B1(n20706), .B2(n2981), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_1/DFF_12/N3 ) );
  AOI22_X1 U20287 ( .A1(n24024), .A2(n26715), .B1(n20632), .B2(n3007), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_13/DFF_12/N3 ) );
  AOI22_X1 U20288 ( .A1(n23997), .A2(n26715), .B1(n20686), .B2(n3003), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_10/DFF_12/N3 ) );
  AOI22_X1 U20289 ( .A1(n24018), .A2(n26715), .B1(n20296), .B2(n2990), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_30/DFF_12/N3 ) );
  AOI22_X1 U20290 ( .A1(n24014), .A2(n26715), .B1(n20668), .B2(n24819), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_11/DFF_12/N3 ) );
  AOI22_X1 U20291 ( .A1(n24011), .A2(n26715), .B1(n20433), .B2(n24825), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_22/DFF_12/N3 ) );
  AOI22_X1 U20292 ( .A1(n24015), .A2(n26715), .B1(n20204), .B2(n3000), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_6/DFF_12/N3 ) );
  AOI22_X1 U20293 ( .A1(n24016), .A2(n26715), .B1(n3001), .B2(n20223), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_5/DFF_12/N3 ) );
  AOI22_X1 U20294 ( .A1(n24002), .A2(n26715), .B1(n20394), .B2(n2988), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_24/DFF_12/N3 ) );
  AOI22_X1 U20295 ( .A1(n23996), .A2(n26715), .B1(n20502), .B2(n2982), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_19/DFF_12/N3 ) );
  AOI22_X1 U20296 ( .A1(n24004), .A2(n26715), .B1(n20351), .B2(n24827), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_28/DFF_12/N3 ) );
  AOI22_X1 U20297 ( .A1(n24005), .A2(n26715), .B1(n20368), .B2(n24620), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_27/DFF_12/N3 ) );
  AOI22_X1 U20298 ( .A1(n23999), .A2(n26715), .B1(n20549), .B2(n24820), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_17/DFF_12/N3 ) );
  AOI22_X1 U20299 ( .A1(n24017), .A2(n26715), .B1(n2997), .B2(n20243), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_4/DFF_12/N3 ) );
  AOI22_X1 U20300 ( .A1(n24022), .A2(n26715), .B1(n20613), .B2(n3006), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_14/DFF_12/N3 ) );
  AOI22_X1 U20301 ( .A1(n24019), .A2(n26715), .B1(n2998), .B2(n20315), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_3/DFF_12/N3 ) );
  AOI22_X1 U20302 ( .A1(n24003), .A2(n26715), .B1(n20375), .B2(n2987), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_25/DFF_12/N3 ) );
  AOI22_X1 U20303 ( .A1(n24020), .A2(n26715), .B1(n20464), .B2(n2985), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_20/DFF_12/N3 ) );
  AOI22_X1 U20304 ( .A1(n24021), .A2(n26715), .B1(n20483), .B2(n2991), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_2/DFF_12/N3 ) );
  AOI22_X1 U20305 ( .A1(n24001), .A2(n26715), .B1(n20445), .B2(n2984), .ZN(
        \core_inst/ID/REGISTER_FILE/REG_21/DFF_12/N3 ) );
  NOR2_X1 U20306 ( .A1(net716333), .A2(n22677), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_26/N3 ) );
  NOR2_X1 U20307 ( .A1(net796193), .A2(n26740), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_0/N3 ) );
  NOR2_X1 U20308 ( .A1(net796114), .A2(net712378), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_5/N3 ) );
  NOR2_X1 U20309 ( .A1(net716313), .A2(n26725), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_3/N3 ) );
  NOR2_X1 U20310 ( .A1(net716311), .A2(n753), .ZN(
        \core_inst/IDEX_NPC/DFF_21/N3 ) );
  NOR2_X1 U20311 ( .A1(net804641), .A2(n26738), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_11/N3 ) );
  NOR2_X1 U20312 ( .A1(net716333), .A2(net712377), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_7/N3 ) );
  NOR2_X1 U20313 ( .A1(net796193), .A2(n26739), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_10/N3 ) );
  OAI211_X1 U20314 ( .C1(n19338), .C2(n624), .A(n26330), .B(n19645), .ZN(
        n26331) );
  NAND2_X1 U20315 ( .A1(n25674), .A2(n24796), .ZN(n26330) );
  NAND2_X1 U20316 ( .A1(n25674), .A2(n24729), .ZN(n26325) );
  NAND2_X1 U20317 ( .A1(n26602), .A2(n26601), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_13/N3 ) );
  AOI211_X1 U20318 ( .C1(n18529), .C2(n997), .A(n26595), .B(n19090), .ZN(
        n26596) );
  OAI22_X1 U20319 ( .A1(n18387), .A2(n2965), .B1(n18400), .B2(n2962), .ZN(
        n26595) );
  NOR2_X1 U20320 ( .A1(n26594), .A2(n26593), .ZN(n26597) );
  OAI211_X1 U20321 ( .C1(n18390), .C2(n2961), .A(n19110), .B(n26592), .ZN(
        n26593) );
  NAND2_X1 U20322 ( .A1(n17796), .A2(net712520), .ZN(n26592) );
  NAND4_X1 U20323 ( .A1(n19107), .A2(n19104), .A3(n19105), .A4(n19106), .ZN(
        n26594) );
  NOR3_X1 U20324 ( .A1(n19093), .A2(n19092), .A3(n19091), .ZN(n26598) );
  OAI21_X1 U20325 ( .B1(n25546), .B2(n25547), .A(n26704), .ZN(n25544) );
  NAND4_X1 U20326 ( .A1(n19916), .A2(n24834), .A3(n19917), .A4(n25548), .ZN(
        n25547) );
  NAND2_X1 U20327 ( .A1(n26663), .A2(n17728), .ZN(n25719) );
  AOI22_X1 U20328 ( .A1(net741608), .A2(n24605), .B1(net712606), .B2(n600), 
        .ZN(n25720) );
  OAI21_X1 U20329 ( .B1(n25538), .B2(n25539), .A(net717052), .ZN(n25536) );
  NAND4_X1 U20330 ( .A1(n25540), .A2(n18725), .A3(n18717), .A4(n18724), .ZN(
        n25539) );
  NOR2_X1 U20331 ( .A1(n25541), .A2(n25542), .ZN(n25540) );
  NOR2_X1 U20332 ( .A1(n18332), .A2(n624), .ZN(n25542) );
  OAI21_X1 U20333 ( .B1(n618), .B2(net767169), .A(n18723), .ZN(n25541) );
  NAND4_X1 U20334 ( .A1(n18706), .A2(n24833), .A3(n18707), .A4(n25543), .ZN(
        n25538) );
  NOR2_X1 U20335 ( .A1(net812958), .A2(n1660), .ZN(
        \core_inst/EXMEM_IR/DFF_13/N3 ) );
  NOR2_X1 U20336 ( .A1(net716333), .A2(n953), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_16/N3 ) );
  OAI21_X1 U20337 ( .B1(n26666), .B2(n26665), .A(n26704), .ZN(n26667) );
  NAND4_X1 U20338 ( .A1(n26664), .A2(n19970), .A3(n19971), .A4(n19969), .ZN(
        n26665) );
  NAND2_X1 U20339 ( .A1(net712499), .A2(n26714), .ZN(n26668) );
  NAND2_X1 U20340 ( .A1(n25665), .A2(n26675), .ZN(n26676) );
  OAI21_X1 U20341 ( .B1(n26674), .B2(n26673), .A(n26704), .ZN(n26677) );
  NAND4_X1 U20342 ( .A1(n19403), .A2(n19400), .A3(n19401), .A4(n19402), .ZN(
        n26673) );
  OAI211_X1 U20343 ( .C1(n26785), .C2(n24778), .A(n19409), .B(n19408), .ZN(
        n26674) );
  NAND2_X1 U20344 ( .A1(net717048), .A2(n26624), .ZN(n26625) );
  OAI21_X1 U20345 ( .B1(n26623), .B2(n26622), .A(n26704), .ZN(n26626) );
  NAND4_X1 U20346 ( .A1(n19544), .A2(n19541), .A3(n19542), .A4(n19543), .ZN(
        n26622) );
  OAI211_X1 U20347 ( .C1(n1442), .C2(n26785), .A(n19550), .B(n19549), .ZN(
        n26623) );
  NAND2_X1 U20348 ( .A1(net712397), .A2(n26669), .ZN(n25525) );
  OAI21_X1 U20349 ( .B1(n25526), .B2(n25527), .A(net717052), .ZN(n25524) );
  NAND4_X1 U20350 ( .A1(n25528), .A2(n25529), .A3(n25530), .A4(n25531), .ZN(
        n25526) );
  AOI22_X1 U20351 ( .A1(n18372), .A2(n17999), .B1(net712520), .B2(n24737), 
        .ZN(n25531) );
  AOI22_X1 U20352 ( .A1(net716423), .A2(n17992), .B1(n18373), .B2(n17998), 
        .ZN(n25530) );
  AOI22_X1 U20353 ( .A1(net767214), .A2(n17995), .B1(net767238), .B2(n17989), 
        .ZN(n25529) );
  AOI22_X1 U20354 ( .A1(net767167), .A2(n24596), .B1(net716461), .B2(n24736), 
        .ZN(n25528) );
  NAND2_X1 U20355 ( .A1(net712499), .A2(n26718), .ZN(n25517) );
  OAI21_X1 U20356 ( .B1(n25518), .B2(n25519), .A(n26704), .ZN(n25516) );
  NAND4_X1 U20357 ( .A1(n19472), .A2(n25520), .A3(n19470), .A4(n19469), .ZN(
        n25519) );
  AOI21_X1 U20358 ( .B1(n19336), .B2(n24789), .A(n25521), .ZN(n25520) );
  OAI21_X1 U20359 ( .B1(n25326), .B2(n26785), .A(n19493), .ZN(n25521) );
  NOR2_X1 U20360 ( .A1(n19365), .A2(n2157), .ZN(n25523) );
  OAI222_X1 U20361 ( .A1(n19350), .A2(n2163), .B1(n25678), .B2(n2160), .C1(
        n2159), .C2(n19370), .ZN(n25522) );
  NAND2_X1 U20362 ( .A1(net717048), .A2(n26678), .ZN(n25533) );
  OAI21_X1 U20363 ( .B1(n25534), .B2(n25535), .A(n26704), .ZN(n25532) );
  NAND4_X1 U20364 ( .A1(n19360), .A2(n19357), .A3(n19358), .A4(n19359), .ZN(
        n25535) );
  OAI211_X1 U20365 ( .C1(n26785), .C2(n24779), .A(n19375), .B(n19374), .ZN(
        n25534) );
  OAI21_X1 U20366 ( .B1(n26525), .B2(n26524), .A(n26717), .ZN(n26528) );
  NAND4_X1 U20367 ( .A1(n26523), .A2(n18586), .A3(n18578), .A4(n18585), .ZN(
        n26524) );
  NOR2_X1 U20368 ( .A1(n26522), .A2(n26521), .ZN(n26523) );
  NOR2_X1 U20369 ( .A1(n18332), .A2(n506), .ZN(n26521) );
  OAI21_X1 U20370 ( .B1(n500), .B2(net767169), .A(n18584), .ZN(n26522) );
  NAND4_X1 U20371 ( .A1(n18567), .A2(n24840), .A3(n18568), .A4(n26520), .ZN(
        n26525) );
  NAND2_X1 U20372 ( .A1(n25601), .A2(n17841), .ZN(n25696) );
  AOI22_X1 U20373 ( .A1(net741609), .A2(n25327), .B1(net741527), .B2(n24814), 
        .ZN(n25697) );
  AOI21_X1 U20374 ( .B1(n26701), .B2(n26700), .A(n24008), .ZN(n26703) );
  NOR2_X1 U20375 ( .A1(n26699), .A2(n26698), .ZN(n26700) );
  OAI222_X1 U20376 ( .A1(n18387), .A2(n2929), .B1(n18400), .B2(n2926), .C1(
        n18390), .C2(n2925), .ZN(n26698) );
  AOI22_X1 U20377 ( .A1(n18529), .A2(n24690), .B1(net712520), .B2(n17829), 
        .ZN(n26697) );
  AOI21_X1 U20378 ( .B1(n26298), .B2(n26297), .A(n24008), .ZN(n26301) );
  NOR2_X1 U20379 ( .A1(n26296), .A2(n26295), .ZN(n26297) );
  OAI222_X1 U20380 ( .A1(n18387), .A2(n3037), .B1(n18400), .B2(n3034), .C1(
        n18390), .C2(n3033), .ZN(n26295) );
  AOI22_X1 U20381 ( .A1(n18529), .A2(n24685), .B1(net712520), .B2(n17863), 
        .ZN(n26294) );
  NOR2_X1 U20382 ( .A1(n26293), .A2(n26292), .ZN(n26298) );
  NOR4_X1 U20383 ( .A1(n26357), .A2(n26356), .A3(n26355), .A4(n26354), .ZN(
        n26358) );
  OAI211_X1 U20384 ( .C1(n19338), .C2(n585), .A(n26353), .B(n19623), .ZN(
        n26356) );
  NAND2_X1 U20385 ( .A1(n19393), .A2(n24797), .ZN(n26353) );
  AOI21_X1 U20386 ( .B1(n26381), .B2(n26380), .A(n24008), .ZN(n26382) );
  NOR2_X1 U20387 ( .A1(n26379), .A2(n26378), .ZN(n26380) );
  OAI222_X1 U20388 ( .A1(n18387), .A2(n3073), .B1(n18400), .B2(n3070), .C1(
        n18390), .C2(n3069), .ZN(n26378) );
  AOI22_X1 U20389 ( .A1(n18529), .A2(n24688), .B1(net712520), .B2(n17880), 
        .ZN(n26377) );
  NOR2_X1 U20390 ( .A1(n26376), .A2(n26375), .ZN(n26381) );
  NOR2_X1 U20391 ( .A1(n26637), .A2(n26399), .ZN(n26402) );
  NOR4_X1 U20392 ( .A1(n26398), .A2(n26397), .A3(n26396), .A4(n26395), .ZN(
        n26399) );
  OAI211_X1 U20393 ( .C1(n19338), .C2(n703), .A(n26394), .B(n19865), .ZN(
        n26397) );
  NAND2_X1 U20394 ( .A1(n19393), .A2(n24730), .ZN(n26394) );
  NOR2_X1 U20395 ( .A1(n26637), .A2(n26427), .ZN(n26429) );
  NOR4_X1 U20396 ( .A1(n26426), .A2(n26425), .A3(n26424), .A4(n26423), .ZN(
        n26427) );
  OAI211_X1 U20397 ( .C1(n19338), .C2(n897), .A(n26422), .B(n19821), .ZN(
        n26425) );
  NAND2_X1 U20398 ( .A1(n25674), .A2(n24731), .ZN(n26422) );
  NOR3_X1 U20399 ( .A1(n26446), .A2(n26445), .A3(n26444), .ZN(n26447) );
  NAND4_X1 U20400 ( .A1(n26443), .A2(n26442), .A3(n20085), .A4(n20092), .ZN(
        n26445) );
  OAI22_X1 U20401 ( .A1(n19385), .A2(n3117), .B1(n26785), .B2(n25263), .ZN(
        n26441) );
  AOI21_X1 U20402 ( .B1(n19530), .B2(n24686), .A(n26440), .ZN(n26443) );
  OAI22_X1 U20403 ( .A1(n19383), .A2(n3125), .B1(n19395), .B2(n3118), .ZN(
        n26440) );
  NOR2_X1 U20404 ( .A1(n26637), .A2(n26389), .ZN(n26391) );
  NOR4_X1 U20405 ( .A1(n26388), .A2(n26387), .A3(n26386), .A4(n26385), .ZN(
        n26389) );
  OAI211_X1 U20406 ( .C1(n546), .C2(n19338), .A(n26384), .B(n19601), .ZN(
        n26387) );
  NAND2_X1 U20407 ( .A1(n25674), .A2(n24799), .ZN(n26384) );
  NAND2_X1 U20408 ( .A1(n25601), .A2(n18036), .ZN(n25686) );
  AOI22_X1 U20409 ( .A1(net741609), .A2(n24781), .B1(net741527), .B2(n24587), 
        .ZN(n25687) );
  AOI21_X1 U20410 ( .B1(n26320), .B2(n26319), .A(n24008), .ZN(n26322) );
  NOR2_X1 U20411 ( .A1(n26318), .A2(n26317), .ZN(n26319) );
  OAI222_X1 U20412 ( .A1(n18387), .A2(n3125), .B1(n18400), .B2(n3118), .C1(
        n18390), .C2(n3117), .ZN(n26317) );
  AOI22_X1 U20413 ( .A1(n18529), .A2(n24686), .B1(net712520), .B2(n18024), 
        .ZN(n26316) );
  NOR2_X1 U20414 ( .A1(n26315), .A2(n26314), .ZN(n26320) );
  NAND2_X1 U20415 ( .A1(net717049), .A2(n26675), .ZN(n26544) );
  NAND2_X1 U20416 ( .A1(n25601), .A2(n17923), .ZN(n25739) );
  AOI22_X1 U20417 ( .A1(net741609), .A2(net365821), .B1(net741527), .B2(
        net366191), .ZN(n25740) );
  OAI21_X1 U20418 ( .B1(n26543), .B2(n26542), .A(n25664), .ZN(n26545) );
  NAND2_X1 U20419 ( .A1(n26541), .A2(n26540), .ZN(n26542) );
  NOR4_X1 U20420 ( .A1(n18425), .A2(n18424), .A3(n18433), .A4(n18410), .ZN(
        n26540) );
  NOR4_X1 U20421 ( .A1(n26539), .A2(n18412), .A3(n18411), .A4(n18413), .ZN(
        n26541) );
  NOR2_X1 U20422 ( .A1(net767172), .A2(n2054), .ZN(n26539) );
  NAND4_X1 U20423 ( .A1(n26538), .A2(n26537), .A3(n26536), .A4(n26535), .ZN(
        n26543) );
  AOI22_X1 U20424 ( .A1(n18372), .A2(n17919), .B1(net712520), .B2(n14399), 
        .ZN(n26535) );
  AOI22_X1 U20425 ( .A1(net716423), .A2(n17912), .B1(n18373), .B2(n17918), 
        .ZN(n26536) );
  AOI22_X1 U20426 ( .A1(net767214), .A2(n17915), .B1(n18398), .B2(n17909), 
        .ZN(n26537) );
  AOI22_X1 U20427 ( .A1(net767167), .A2(n24726), .B1(net716461), .B2(n24600), 
        .ZN(n26538) );
  NAND2_X1 U20428 ( .A1(net712397), .A2(n26624), .ZN(n26372) );
  NAND2_X1 U20429 ( .A1(n25601), .A2(n17987), .ZN(n25727) );
  AOI22_X1 U20430 ( .A1(net741609), .A2(net741329), .B1(net741527), .B2(n5307), 
        .ZN(n25728) );
  OAI21_X1 U20431 ( .B1(n26371), .B2(n26370), .A(net717052), .ZN(n26373) );
  NAND2_X1 U20432 ( .A1(n26369), .A2(n26368), .ZN(n26370) );
  NOR4_X1 U20433 ( .A1(n18610), .A2(n18609), .A3(n18618), .A4(n18596), .ZN(
        n26368) );
  NOR4_X1 U20434 ( .A1(n26367), .A2(n18598), .A3(n18597), .A4(n18599), .ZN(
        n26369) );
  NOR2_X1 U20435 ( .A1(net767172), .A2(n2198), .ZN(n26367) );
  NAND4_X1 U20436 ( .A1(n26366), .A2(n26365), .A3(n26364), .A4(n26363), .ZN(
        n26371) );
  AOI22_X1 U20437 ( .A1(n18372), .A2(n17983), .B1(net712520), .B2(n24805), 
        .ZN(n26363) );
  AOI22_X1 U20438 ( .A1(net716423), .A2(n17976), .B1(n18373), .B2(n17982), 
        .ZN(n26364) );
  AOI22_X1 U20439 ( .A1(net767214), .A2(n17979), .B1(n18398), .B2(n17973), 
        .ZN(n26365) );
  AOI22_X1 U20440 ( .A1(net767167), .A2(n24725), .B1(net716461), .B2(n24599), 
        .ZN(n26366) );
  NAND2_X1 U20441 ( .A1(net712499), .A2(n26600), .ZN(n26289) );
  NAND2_X1 U20442 ( .A1(n25601), .A2(n17807), .ZN(n25694) );
  AOI22_X1 U20443 ( .A1(net741609), .A2(n24782), .B1(net741527), .B2(n991), 
        .ZN(n25695) );
  NAND2_X1 U20444 ( .A1(n26704), .A2(n26288), .ZN(n26290) );
  AOI211_X1 U20445 ( .C1(n19530), .C2(n997), .A(n19937), .B(n26284), .ZN(
        n26285) );
  OAI22_X1 U20446 ( .A1(n19383), .A2(n2965), .B1(n19395), .B2(n2962), .ZN(
        n26284) );
  NOR3_X1 U20447 ( .A1(n19940), .A2(n19938), .A3(n19939), .ZN(n26286) );
  AOI211_X1 U20448 ( .C1(n19328), .C2(n24794), .A(n26283), .B(n26282), .ZN(
        n26287) );
  NAND4_X1 U20449 ( .A1(n19950), .A2(n19947), .A3(n19948), .A4(n19949), .ZN(
        n26282) );
  OAI21_X1 U20450 ( .B1(n26785), .B2(n25305), .A(n19952), .ZN(n26283) );
  NAND2_X1 U20451 ( .A1(n25665), .A2(n26669), .ZN(n26620) );
  NAND2_X1 U20452 ( .A1(n26663), .A2(n18003), .ZN(n25708) );
  OAI21_X1 U20453 ( .B1(n26619), .B2(n26618), .A(n26704), .ZN(n26621) );
  NAND2_X1 U20454 ( .A1(n26617), .A2(n26616), .ZN(n26618) );
  NOR4_X1 U20455 ( .A1(n19794), .A2(n19793), .A3(n19801), .A4(n19787), .ZN(
        n26616) );
  NOR4_X1 U20456 ( .A1(n26615), .A2(n19789), .A3(n19788), .A4(n19790), .ZN(
        n26617) );
  NOR2_X1 U20457 ( .A1(n26614), .A2(n2306), .ZN(n26615) );
  NAND4_X1 U20458 ( .A1(n26613), .A2(n26612), .A3(n26611), .A4(n26610), .ZN(
        n26619) );
  AOI22_X1 U20459 ( .A1(n19372), .A2(n17999), .B1(n26609), .B2(n24737), .ZN(
        n26610) );
  AOI22_X1 U20460 ( .A1(n24007), .A2(n17992), .B1(n17998), .B2(n19373), .ZN(
        n26611) );
  AOI22_X1 U20461 ( .A1(n25681), .A2(n17995), .B1(n17989), .B2(n25674), .ZN(
        n26612) );
  AOI22_X1 U20462 ( .A1(n19332), .A2(n24596), .B1(n25679), .B2(n24736), .ZN(
        n26613) );
  NAND2_X1 U20463 ( .A1(net717048), .A2(n26555), .ZN(n26556) );
  OAI21_X1 U20464 ( .B1(n26554), .B2(n26553), .A(n26704), .ZN(n26557) );
  NAND2_X1 U20465 ( .A1(n26552), .A2(n26551), .ZN(n26553) );
  NOR4_X1 U20466 ( .A1(n19456), .A2(n19455), .A3(n19463), .A4(n19449), .ZN(
        n26551) );
  NOR4_X1 U20467 ( .A1(n26550), .A2(n19451), .A3(n19450), .A4(n19452), .ZN(
        n26552) );
  NOR2_X1 U20468 ( .A1(n26614), .A2(n2126), .ZN(n26550) );
  NAND4_X1 U20469 ( .A1(n26549), .A2(n26548), .A3(n26547), .A4(n26546), .ZN(
        n26554) );
  AOI22_X1 U20470 ( .A1(n19372), .A2(n17951), .B1(n26609), .B2(n14401), .ZN(
        n26546) );
  AOI22_X1 U20471 ( .A1(n24007), .A2(n17944), .B1(n19373), .B2(n17950), .ZN(
        n26547) );
  AOI22_X1 U20472 ( .A1(n25681), .A2(n17947), .B1(n25674), .B2(n17941), .ZN(
        n26548) );
  AOI22_X1 U20473 ( .A1(n19332), .A2(n24595), .B1(n25679), .B2(n24735), .ZN(
        n26549) );
  NAND2_X1 U20474 ( .A1(net717049), .A2(n26555), .ZN(n26268) );
  NAND2_X1 U20475 ( .A1(n25601), .A2(n17955), .ZN(n25735) );
  AOI22_X1 U20476 ( .A1(net741609), .A2(net365826), .B1(net741527), .B2(
        net366478), .ZN(n25736) );
  OAI21_X1 U20477 ( .B1(n26267), .B2(n26266), .A(n26717), .ZN(n26269) );
  NAND2_X1 U20478 ( .A1(n26265), .A2(n26264), .ZN(n26266) );
  NOR4_X1 U20479 ( .A1(n18489), .A2(n18488), .A3(n18497), .A4(n18474), .ZN(
        n26264) );
  NOR4_X1 U20480 ( .A1(n26263), .A2(n18476), .A3(n18475), .A4(n18477), .ZN(
        n26265) );
  NOR2_X1 U20481 ( .A1(net767172), .A2(n2126), .ZN(n26263) );
  NAND4_X1 U20482 ( .A1(n26262), .A2(n26261), .A3(n26260), .A4(n26259), .ZN(
        n26267) );
  AOI22_X1 U20483 ( .A1(n18372), .A2(n17951), .B1(net712520), .B2(n14401), 
        .ZN(n26259) );
  AOI22_X1 U20484 ( .A1(net716423), .A2(n17944), .B1(n18373), .B2(n17950), 
        .ZN(n26260) );
  AOI22_X1 U20485 ( .A1(net767214), .A2(n17947), .B1(net767238), .B2(n17941), 
        .ZN(n26261) );
  AOI22_X1 U20486 ( .A1(net767167), .A2(n24595), .B1(net716461), .B2(n24735), 
        .ZN(n26262) );
  NAND2_X1 U20487 ( .A1(n25665), .A2(n26639), .ZN(n26503) );
  NAND2_X1 U20488 ( .A1(n25601), .A2(n17939), .ZN(n25737) );
  AOI22_X1 U20489 ( .A1(net741609), .A2(n24780), .B1(net741527), .B2(n5729), 
        .ZN(n25738) );
  OAI21_X1 U20490 ( .B1(n26502), .B2(n26501), .A(n26704), .ZN(n26504) );
  NAND2_X1 U20491 ( .A1(n26500), .A2(n26499), .ZN(n26501) );
  NOR4_X1 U20492 ( .A1(n19434), .A2(n19433), .A3(n19441), .A4(n19427), .ZN(
        n26499) );
  NOR4_X1 U20493 ( .A1(n26498), .A2(n19429), .A3(n19428), .A4(n19430), .ZN(
        n26500) );
  NOR2_X1 U20494 ( .A1(n26614), .A2(n2090), .ZN(n26498) );
  NAND4_X1 U20495 ( .A1(n26497), .A2(n26496), .A3(n26495), .A4(n26494), .ZN(
        n26502) );
  AOI22_X1 U20496 ( .A1(n19372), .A2(n17935), .B1(n26609), .B2(n14127), .ZN(
        n26494) );
  AOI22_X1 U20497 ( .A1(n24007), .A2(n17928), .B1(n17934), .B2(n19373), .ZN(
        n26495) );
  AOI22_X1 U20498 ( .A1(n25681), .A2(n17931), .B1(n17925), .B2(n25674), .ZN(
        n26496) );
  AOI22_X1 U20499 ( .A1(n24026), .A2(n24597), .B1(n25679), .B2(n24738), .ZN(
        n26497) );
  NAND2_X1 U20500 ( .A1(net717050), .A2(n26678), .ZN(n26343) );
  NAND2_X1 U20501 ( .A1(n25601), .A2(n17908), .ZN(n25741) );
  OAI21_X1 U20502 ( .B1(n26342), .B2(n26341), .A(net717052), .ZN(n26344) );
  NAND2_X1 U20503 ( .A1(n26340), .A2(n26339), .ZN(n26341) );
  NOR4_X1 U20504 ( .A1(n18381), .A2(n18380), .A3(n18399), .A4(n18357), .ZN(
        n26339) );
  NOR4_X1 U20505 ( .A1(n26338), .A2(n18359), .A3(n18358), .A4(n18360), .ZN(
        n26340) );
  NOR2_X1 U20506 ( .A1(net767172), .A2(n2018), .ZN(n26338) );
  NAND4_X1 U20507 ( .A1(n26337), .A2(n26336), .A3(n26335), .A4(n26334), .ZN(
        n26342) );
  AOI22_X1 U20508 ( .A1(n18372), .A2(n17904), .B1(net712520), .B2(n14400), 
        .ZN(n26334) );
  AOI22_X1 U20509 ( .A1(net716423), .A2(n17897), .B1(n18373), .B2(n17903), 
        .ZN(n26335) );
  AOI22_X1 U20510 ( .A1(net767214), .A2(n17900), .B1(n18398), .B2(n17894), 
        .ZN(n26336) );
  AOI22_X1 U20511 ( .A1(net767167), .A2(n24724), .B1(net716461), .B2(n24598), 
        .ZN(n26337) );
  NAND2_X1 U20512 ( .A1(n25601), .A2(n17706), .ZN(n25729) );
  AOI22_X1 U20513 ( .A1(net741609), .A2(n25328), .B1(net741527), .B2(n482), 
        .ZN(n25730) );
  NOR2_X1 U20514 ( .A1(n26637), .A2(n26309), .ZN(n26311) );
  NOR4_X1 U20515 ( .A1(n26308), .A2(n26307), .A3(n26306), .A4(n26305), .ZN(
        n26309) );
  OAI211_X1 U20516 ( .C1(n19338), .C2(n506), .A(n26304), .B(n19535), .ZN(
        n26307) );
  NAND2_X1 U20517 ( .A1(n25674), .A2(n24795), .ZN(n26304) );
  NAND2_X1 U20518 ( .A1(n25601), .A2(n17699), .ZN(n25731) );
  AOI22_X1 U20519 ( .A1(net741609), .A2(n24773), .B1(net741527), .B2(net741582), .ZN(n25732) );
  NAND2_X1 U20520 ( .A1(n25674), .A2(n24798), .ZN(n26359) );
  NAND4_X1 U20521 ( .A1(n19500), .A2(n19502), .A3(n19499), .A4(n19501), .ZN(
        n26361) );
  NOR2_X1 U20522 ( .A1(n26680), .A2(n26679), .ZN(n26681) );
  NOR2_X1 U20523 ( .A1(n18332), .A2(n356), .ZN(n26679) );
  OAI21_X1 U20524 ( .B1(n350), .B2(net767169), .A(n18334), .ZN(n26680) );
  NAND4_X1 U20525 ( .A1(n18299), .A2(n18296), .A3(n18297), .A4(n18298), .ZN(
        n26683) );
  AOI21_X1 U20526 ( .B1(n26693), .B2(n26692), .A(n24008), .ZN(n26695) );
  NOR2_X1 U20527 ( .A1(n26691), .A2(n26690), .ZN(n26692) );
  OAI222_X1 U20528 ( .A1(n18387), .A2(n3001), .B1(n18400), .B2(n2998), .C1(
        n18390), .C2(n2997), .ZN(n26690) );
  AOI22_X1 U20529 ( .A1(n18529), .A2(n24681), .B1(net712520), .B2(n17846), 
        .ZN(n26689) );
  NOR2_X1 U20530 ( .A1(n26688), .A2(n26687), .ZN(n26693) );
  NOR2_X1 U20531 ( .A1(n26608), .A2(n26607), .ZN(net712377) );
  AOI21_X1 U20532 ( .B1(n6462), .B2(net712812), .A(n26570), .ZN(n26257) );
  NOR2_X1 U20533 ( .A1(n26637), .A2(n26477), .ZN(n26480) );
  NOR4_X1 U20534 ( .A1(n26476), .A2(n26475), .A3(n26474), .A4(n26473), .ZN(
        n26477) );
  OAI211_X1 U20535 ( .C1(n19338), .C2(n779), .A(n26472), .B(n19711), .ZN(
        n26475) );
  NAND2_X1 U20536 ( .A1(n25674), .A2(n24733), .ZN(n26472) );
  NAND2_X1 U20537 ( .A1(n26663), .A2(n17763), .ZN(net715885) );
  AOI22_X1 U20538 ( .A1(net741608), .A2(n5664), .B1(net712606), .B2(n794), 
        .ZN(net715884) );
  NOR4_X1 U20539 ( .A1(n26454), .A2(n26453), .A3(n26452), .A4(n26451), .ZN(
        n26455) );
  OAI211_X1 U20540 ( .C1(n19338), .C2(n818), .A(n26450), .B(n19733), .ZN(
        n26453) );
  NAND2_X1 U20541 ( .A1(n25674), .A2(net741400), .ZN(n26450) );
  NOR2_X1 U20542 ( .A1(n26637), .A2(n26466), .ZN(n26469) );
  NOR4_X1 U20543 ( .A1(n26465), .A2(n26464), .A3(n26463), .A4(n26462), .ZN(
        n26466) );
  OAI211_X1 U20544 ( .C1(n19338), .C2(n394), .A(n26461), .B(n19667), .ZN(
        n26464) );
  NAND2_X1 U20545 ( .A1(n25674), .A2(n24732), .ZN(n26461) );
  OAI211_X1 U20546 ( .C1(n936), .C2(n19338), .A(n26633), .B(n19843), .ZN(
        n26635) );
  NAND2_X1 U20547 ( .A1(n19393), .A2(n24803), .ZN(n26633) );
  NAND2_X1 U20548 ( .A1(n25601), .A2(n17892), .ZN(n25690) );
  AOI22_X1 U20549 ( .A1(net741609), .A2(n24806), .B1(net741527), .B2(n24601), 
        .ZN(n25691) );
  NOR3_X1 U20550 ( .A1(n26629), .A2(n26628), .A3(n26627), .ZN(n26630) );
  NOR2_X1 U20551 ( .A1(n26637), .A2(n26417), .ZN(n26419) );
  NOR4_X1 U20552 ( .A1(n26416), .A2(n26415), .A3(n26414), .A4(n26413), .ZN(
        n26417) );
  OAI211_X1 U20553 ( .C1(n19338), .C2(n664), .A(n26412), .B(n19689), .ZN(
        n26415) );
  NAND2_X1 U20554 ( .A1(n19393), .A2(n24734), .ZN(n26412) );
  NOR2_X1 U20555 ( .A1(n26637), .A2(n26589), .ZN(n26591) );
  NOR4_X1 U20556 ( .A1(n26588), .A2(n26587), .A3(n26586), .A4(n26585), .ZN(
        n26589) );
  OAI211_X1 U20557 ( .C1(n432), .C2(n19338), .A(n26584), .B(n19579), .ZN(
        n26587) );
  NAND2_X1 U20558 ( .A1(n25674), .A2(n24802), .ZN(n26584) );
  AOI21_X1 U20559 ( .B1(n26489), .B2(n26488), .A(n24008), .ZN(n26492) );
  NOR2_X1 U20560 ( .A1(n26487), .A2(n26486), .ZN(n26488) );
  OAI222_X1 U20561 ( .A1(n18387), .A2(n2713), .B1(n18400), .B2(n2710), .C1(
        n18390), .C2(n2709), .ZN(n26486) );
  AOI22_X1 U20562 ( .A1(n18529), .A2(n24687), .B1(net712520), .B2(n18007), 
        .ZN(n26485) );
  NOR2_X1 U20563 ( .A1(n26484), .A2(n26483), .ZN(n26489) );
  NAND2_X1 U20564 ( .A1(n26663), .A2(n17770), .ZN(n25709) );
  AOI22_X1 U20565 ( .A1(net741608), .A2(n24808), .B1(net712606), .B2(n834), 
        .ZN(n25710) );
  NOR2_X1 U20566 ( .A1(n26637), .A2(n26517), .ZN(n26518) );
  NOR4_X1 U20567 ( .A1(n26516), .A2(n26515), .A3(n26514), .A4(n26513), .ZN(
        n26517) );
  OAI211_X1 U20568 ( .C1(n19338), .C2(n858), .A(n26512), .B(n19777), .ZN(
        n26515) );
  NAND2_X1 U20569 ( .A1(n25674), .A2(net741397), .ZN(n26512) );
  NAND2_X1 U20570 ( .A1(n25601), .A2(n17824), .ZN(n25698) );
  AOI22_X1 U20571 ( .A1(net741609), .A2(n24606), .B1(net741527), .B2(n24810), 
        .ZN(n25699) );
  AOI21_X1 U20572 ( .B1(n26647), .B2(n26646), .A(n24008), .ZN(n26650) );
  NOR2_X1 U20573 ( .A1(n26645), .A2(n26644), .ZN(n26646) );
  OAI222_X1 U20574 ( .A1(n18387), .A2(n2893), .B1(n18400), .B2(n2890), .C1(
        n18390), .C2(n2889), .ZN(n26644) );
  AOI22_X1 U20575 ( .A1(n18529), .A2(n24689), .B1(net712520), .B2(n17812), 
        .ZN(n26643) );
  NOR2_X1 U20576 ( .A1(n26642), .A2(n26641), .ZN(n26647) );
  NAND2_X1 U20577 ( .A1(n25601), .A2(n17682), .ZN(n25742) );
  AOI22_X1 U20578 ( .A1(net741609), .A2(n24809), .B1(net741527), .B2(n5761), 
        .ZN(n25743) );
  NOR2_X1 U20579 ( .A1(n26637), .A2(n26505), .ZN(n26507) );
  NAND2_X1 U20580 ( .A1(n26663), .A2(n17750), .ZN(n25711) );
  AOI22_X1 U20581 ( .A1(net741608), .A2(n25329), .B1(net712606), .B2(n717), 
        .ZN(n25712) );
  OAI21_X1 U20582 ( .B1(n25559), .B2(n25560), .A(n25664), .ZN(n25557) );
  NAND4_X1 U20583 ( .A1(n25561), .A2(n18860), .A3(n18852), .A4(n18859), .ZN(
        n25560) );
  NOR2_X1 U20584 ( .A1(n25562), .A2(n25563), .ZN(n25561) );
  NOR2_X1 U20585 ( .A1(n18332), .A2(n741), .ZN(n25563) );
  OAI21_X1 U20586 ( .B1(n735), .B2(net767169), .A(n18858), .ZN(n25562) );
  NAND4_X1 U20587 ( .A1(n18841), .A2(n24836), .A3(n18842), .A4(n25564), .ZN(
        n25559) );
  NAND2_X1 U20588 ( .A1(n26663), .A2(n17784), .ZN(n25704) );
  AOI22_X1 U20589 ( .A1(net741608), .A2(n25330), .B1(net712606), .B2(n912), 
        .ZN(n25705) );
  OAI21_X1 U20590 ( .B1(n25571), .B2(n25572), .A(n25664), .ZN(n25569) );
  NAND4_X1 U20591 ( .A1(n25573), .A2(n18972), .A3(n18964), .A4(n18971), .ZN(
        n25572) );
  NOR2_X1 U20592 ( .A1(n25574), .A2(n25575), .ZN(n25573) );
  NOR2_X1 U20593 ( .A1(n18332), .A2(n936), .ZN(n25575) );
  OAI21_X1 U20594 ( .B1(n930), .B2(net767169), .A(n18970), .ZN(n25574) );
  NAND2_X1 U20595 ( .A1(n26663), .A2(n17695), .ZN(n25725) );
  AOI22_X1 U20596 ( .A1(net741608), .A2(n24604), .B1(net712606), .B2(n24817), 
        .ZN(n25726) );
  OAI21_X1 U20597 ( .B1(n25551), .B2(n25552), .A(n25664), .ZN(n25549) );
  NAND4_X1 U20598 ( .A1(n25553), .A2(n18644), .A3(n18636), .A4(n18643), .ZN(
        n25552) );
  NOR2_X1 U20599 ( .A1(n25554), .A2(n25555), .ZN(n25553) );
  NOR2_X1 U20600 ( .A1(n18332), .A2(n432), .ZN(n25555) );
  OAI21_X1 U20601 ( .B1(n426), .B2(net767169), .A(n18642), .ZN(n25554) );
  NAND4_X1 U20602 ( .A1(n18625), .A2(n24835), .A3(n18626), .A4(n25556), .ZN(
        n25551) );
  NAND2_X1 U20603 ( .A1(n25601), .A2(n17971), .ZN(n25733) );
  AOI22_X1 U20604 ( .A1(net741609), .A2(n24602), .B1(net741527), .B2(net741305), .ZN(n25734) );
  OAI21_X1 U20605 ( .B1(n25567), .B2(n25568), .A(net717052), .ZN(n25565) );
  NOR2_X1 U20606 ( .A1(net812952), .A2(net712353), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_12/N3 ) );
  INV_X1 U20607 ( .A(net712445), .ZN(net712353) );
  NOR2_X1 U20608 ( .A1(net716313), .A2(n24787), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_27/N3 ) );
  NOR2_X1 U20609 ( .A1(net716333), .A2(net712356), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_25/N3 ) );
  NAND2_X1 U20610 ( .A1(n26663), .A2(n17735), .ZN(n25715) );
  AOI22_X1 U20611 ( .A1(net741608), .A2(n25337), .B1(net712606), .B2(n640), 
        .ZN(n25716) );
  OAI21_X1 U20612 ( .B1(n26657), .B2(n26656), .A(n26717), .ZN(n26660) );
  NAND4_X1 U20613 ( .A1(n25262), .A2(n18779), .A3(n18771), .A4(n18778), .ZN(
        n26656) );
  NAND2_X1 U20614 ( .A1(net767238), .A2(n24734), .ZN(n26654) );
  NAND4_X1 U20615 ( .A1(n18760), .A2(n24841), .A3(n18761), .A4(n26653), .ZN(
        n26657) );
  NAND2_X1 U20616 ( .A1(n25601), .A2(n17742), .ZN(n25702) );
  AOI22_X1 U20617 ( .A1(net741609), .A2(n25317), .B1(net741527), .B2(n679), 
        .ZN(n25703) );
  OAI21_X1 U20618 ( .B1(n26349), .B2(n26348), .A(n26717), .ZN(n26351) );
  NAND4_X1 U20619 ( .A1(n25261), .A2(n18999), .A3(n18991), .A4(n18998), .ZN(
        n26348) );
  NAND2_X1 U20620 ( .A1(n18398), .A2(n24730), .ZN(n26346) );
  NAND4_X1 U20621 ( .A1(n18980), .A2(n24838), .A3(n18981), .A4(n26345), .ZN(
        n26349) );
  NAND2_X1 U20622 ( .A1(n26663), .A2(n17720), .ZN(n25721) );
  AOI22_X1 U20623 ( .A1(net741608), .A2(n24783), .B1(net712606), .B2(n561), 
        .ZN(n25722) );
  OAI21_X1 U20624 ( .B1(n26435), .B2(n26434), .A(n25664), .ZN(n26438) );
  NAND4_X1 U20625 ( .A1(n26433), .A2(n18698), .A3(n18690), .A4(n18697), .ZN(
        n26434) );
  NOR2_X1 U20626 ( .A1(n26432), .A2(n26431), .ZN(n26433) );
  NOR2_X1 U20627 ( .A1(n18332), .A2(n585), .ZN(n26431) );
  OAI21_X1 U20628 ( .B1(n579), .B2(net767169), .A(n18696), .ZN(n26432) );
  NAND4_X1 U20629 ( .A1(n18679), .A2(n24839), .A3(n18680), .A4(n26430), .ZN(
        n26435) );
  NAND2_X1 U20630 ( .A1(n26663), .A2(n17688), .ZN(n25717) );
  AOI22_X1 U20631 ( .A1(net741608), .A2(n24603), .B1(net712606), .B2(n24816), 
        .ZN(n25718) );
  NAND2_X1 U20632 ( .A1(n26663), .A2(n17713), .ZN(n25723) );
  AOI22_X1 U20633 ( .A1(net741608), .A2(n24784), .B1(net712606), .B2(n522), 
        .ZN(n25724) );
  NAND2_X1 U20634 ( .A1(n26663), .A2(n17777), .ZN(n25706) );
  AOI22_X1 U20635 ( .A1(net741608), .A2(net741301), .B1(net712606), .B2(n873), 
        .ZN(n25707) );
  NAND2_X1 U20636 ( .A1(n26663), .A2(n17756), .ZN(n25713) );
  AOI22_X1 U20637 ( .A1(net741608), .A2(n25318), .B1(net712606), .B2(n755), 
        .ZN(n25714) );
  OAI21_X1 U20638 ( .B1(n26279), .B2(n26278), .A(n25664), .ZN(n26281) );
  NAND4_X1 U20639 ( .A1(n25260), .A2(n18806), .A3(n18798), .A4(n18805), .ZN(
        n26278) );
  NAND2_X1 U20640 ( .A1(net767238), .A2(n24733), .ZN(n26276) );
  NAND4_X1 U20641 ( .A1(n18787), .A2(n24837), .A3(n18788), .A4(n26275), .ZN(
        n26279) );
  NAND2_X1 U20642 ( .A1(n25601), .A2(n18019), .ZN(n25688) );
  AOI22_X1 U20643 ( .A1(net741609), .A2(n25319), .B1(net741527), .B2(net366126), .ZN(n25689) );
  NAND2_X1 U20644 ( .A1(n25601), .A2(n17791), .ZN(n25700) );
  AOI22_X1 U20645 ( .A1(net741609), .A2(n24807), .B1(net741527), .B2(n952), 
        .ZN(n25701) );
  NAND2_X1 U20646 ( .A1(n25601), .A2(n17875), .ZN(n25692) );
  AOI22_X1 U20647 ( .A1(net741609), .A2(n24607), .B1(net741527), .B2(n24812), 
        .ZN(n25693) );
  NAND2_X1 U20648 ( .A1(n20061), .A2(n20077), .ZN(n19385) );
  NAND2_X1 U20649 ( .A1(n26776), .A2(s_IFID_IR[26]), .ZN(net518455) );
  NOR2_X1 U20650 ( .A1(net716311), .A2(n26737), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_17/N3 ) );
  NAND2_X1 U20651 ( .A1(s_IFID_IR[30]), .A2(n19282), .ZN(n20118) );
  NAND2_X1 U20652 ( .A1(n18133), .A2(n18132), .ZN(net712961) );
  NAND2_X1 U20653 ( .A1(n25745), .A2(n18175), .ZN(n18135) );
  NAND2_X1 U20654 ( .A1(n24584), .A2(n24813), .ZN(n26511) );
  NOR2_X1 U20655 ( .A1(s_IFID_IR[26]), .A2(n18171), .ZN(n26258) );
  OAI21_X1 U20656 ( .B1(net741531), .B2(net366211), .A(net716215), .ZN(n26255)
         );
  NOR3_X1 U20657 ( .A1(n26233), .A2(net713554), .A3(net713151), .ZN(n26239) );
  NAND2_X1 U20658 ( .A1(n24358), .A2(n23975), .ZN(n26215) );
  NAND2_X1 U20659 ( .A1(n24274), .A2(n24318), .ZN(n26187) );
  NAND2_X1 U20660 ( .A1(net713767), .A2(n26169), .ZN(n26170) );
  NOR2_X1 U20661 ( .A1(n26168), .A2(net713770), .ZN(n26171) );
  NAND2_X1 U20662 ( .A1(net718367), .A2(net713775), .ZN(n26166) );
  AOI22_X1 U20663 ( .A1(n26153), .A2(n26152), .B1(n24306), .B2(n23975), .ZN(
        n26164) );
  NAND2_X1 U20664 ( .A1(net713829), .A2(net713151), .ZN(n26405) );
  NOR2_X1 U20665 ( .A1(net713905), .A2(n26133), .ZN(net713930) );
  AOI21_X1 U20666 ( .B1(net712466), .B2(net749685), .A(n25406), .ZN(n26124) );
  NOR2_X1 U20667 ( .A1(n26122), .A2(n26121), .ZN(n26125) );
  NOR4_X1 U20668 ( .A1(n26114), .A2(n26113), .A3(n22800), .A4(n26111), .ZN(
        n26115) );
  NOR4_X1 U20669 ( .A1(n26109), .A2(n26108), .A3(n26107), .A4(n26106), .ZN(
        n26116) );
  NOR2_X1 U20670 ( .A1(n26104), .A2(n26103), .ZN(n26117) );
  NAND4_X1 U20671 ( .A1(n24325), .A2(n26102), .A3(n24087), .A4(n24289), .ZN(
        n26103) );
  NOR3_X1 U20672 ( .A1(n26092), .A2(n24553), .A3(n26091), .ZN(n26093) );
  NOR4_X1 U20673 ( .A1(n26087), .A2(n26086), .A3(n26085), .A4(n26084), .ZN(
        n26094) );
  NOR2_X1 U20674 ( .A1(n26083), .A2(n26082), .ZN(n26095) );
  NAND4_X1 U20675 ( .A1(n26081), .A2(net742296), .A3(net749295), .A4(net762762), .ZN(n26082) );
  NAND2_X1 U20676 ( .A1(n25476), .A2(n25477), .ZN(n25475) );
  OAI22_X1 U20677 ( .A1(net714182), .A2(n24328), .B1(n26066), .B2(net767210), 
        .ZN(n25473) );
  NOR3_X1 U20678 ( .A1(n25478), .A2(n25479), .A3(n25480), .ZN(net714174) );
  NOR3_X1 U20679 ( .A1(net749812), .A2(n24357), .A3(net767203), .ZN(n25480) );
  NAND4_X1 U20680 ( .A1(n25481), .A2(n25482), .A3(n25483), .A4(n25484), .ZN(
        n25478) );
  NAND4_X1 U20681 ( .A1(n25490), .A2(n25491), .A3(n25492), .A4(n25493), .ZN(
        n25485) );
  NAND2_X1 U20682 ( .A1(n24312), .A2(net713736), .ZN(n25495) );
  NAND2_X1 U20683 ( .A1(n26060), .A2(net713892), .ZN(n25494) );
  NAND2_X1 U20684 ( .A1(n26059), .A2(n26056), .ZN(n25491) );
  AOI22_X1 U20685 ( .A1(n26136), .A2(n26190), .B1(n26214), .B2(net767234), 
        .ZN(n25490) );
  NAND2_X1 U20686 ( .A1(n26056), .A2(net718367), .ZN(n25376) );
  NAND2_X1 U20687 ( .A1(n25468), .A2(net750032), .ZN(n25500) );
  NOR2_X1 U20688 ( .A1(n24546), .A2(net767203), .ZN(n25468) );
  XNOR2_X1 U20689 ( .A(n24178), .B(n24274), .ZN(n26037) );
  NOR2_X1 U20690 ( .A1(n26014), .A2(n26013), .ZN(n26017) );
  OAI21_X1 U20691 ( .B1(net366531), .B2(net713775), .A(n26012), .ZN(n26013) );
  NOR2_X1 U20692 ( .A1(n25467), .A2(n26008), .ZN(n25445) );
  NAND2_X1 U20693 ( .A1(n26163), .A2(net767211), .ZN(n26015) );
  NAND2_X1 U20694 ( .A1(n26050), .A2(net713785), .ZN(n26011) );
  NOR4_X1 U20695 ( .A1(n26010), .A2(n26006), .A3(n26005), .A4(n26004), .ZN(
        n26007) );
  NOR2_X1 U20696 ( .A1(n26031), .A2(net755699), .ZN(n26005) );
  OAI22_X1 U20697 ( .A1(net713810), .A2(net796212), .B1(n24357), .B2(net713773), .ZN(n26006) );
  NAND2_X1 U20698 ( .A1(n25965), .A2(n25964), .ZN(n26533) );
  NOR2_X1 U20699 ( .A1(n25963), .A2(n25962), .ZN(n25964) );
  NOR2_X1 U20700 ( .A1(n23974), .A2(net713726), .ZN(n25961) );
  OAI22_X1 U20701 ( .A1(net714261), .A2(net713897), .B1(net713738), .B2(n26196), .ZN(n25963) );
  NOR2_X1 U20702 ( .A1(n25938), .A2(n22871), .ZN(n25503) );
  AOI21_X1 U20703 ( .B1(n25883), .B2(n25882), .A(net767203), .ZN(n25895) );
  NOR3_X1 U20704 ( .A1(n25879), .A2(n25878), .A3(n25877), .ZN(n25883) );
  NAND2_X1 U20705 ( .A1(n26041), .A2(n24313), .ZN(n25876) );
  NOR3_X1 U20706 ( .A1(n25930), .A2(n25929), .A3(n25928), .ZN(n25931) );
  NOR3_X1 U20707 ( .A1(n25927), .A2(n25926), .A3(n25925), .ZN(n25932) );
  OAI21_X1 U20708 ( .B1(n25924), .B2(net714476), .A(n25923), .ZN(n25927) );
  AOI21_X1 U20709 ( .B1(n25917), .B2(n25916), .A(net767203), .ZN(n25918) );
  NOR3_X1 U20710 ( .A1(n25915), .A2(n25914), .A3(n25913), .ZN(n25916) );
  NOR3_X1 U20711 ( .A1(n25912), .A2(n25911), .A3(n25910), .ZN(n25917) );
  OAI22_X1 U20712 ( .A1(n24177), .A2(net767210), .B1(n26066), .B2(net714182), 
        .ZN(n25902) );
  NOR2_X1 U20713 ( .A1(n25874), .A2(n24097), .ZN(n26560) );
  AOI21_X1 U20714 ( .B1(n26127), .B2(n25873), .A(n26129), .ZN(n26566) );
  NAND2_X1 U20715 ( .A1(n25381), .A2(n25865), .ZN(n25867) );
  NAND2_X1 U20716 ( .A1(n26218), .A2(n24173), .ZN(n25862) );
  XNOR2_X1 U20717 ( .A(n22696), .B(net713564), .ZN(net714335) );
  NOR2_X1 U20718 ( .A1(n24353), .A2(n26118), .ZN(n25472) );
  NAND4_X1 U20719 ( .A1(n25820), .A2(n25819), .A3(n25818), .A4(n25817), .ZN(
        n26607) );
  AOI22_X1 U20720 ( .A1(n24545), .A2(net714306), .B1(net767234), .B2(n26186), 
        .ZN(n25818) );
  AOI21_X1 U20721 ( .B1(n25814), .B2(net713775), .A(n25813), .ZN(n25820) );
  NAND2_X1 U20722 ( .A1(n25381), .A2(n25810), .ZN(n25811) );
  NOR2_X1 U20723 ( .A1(n24531), .A2(net717087), .ZN(n25812) );
  NAND4_X1 U20724 ( .A1(n25809), .A2(n25808), .A3(n25807), .A4(n25806), .ZN(
        n25814) );
  NAND2_X1 U20725 ( .A1(n25596), .A2(net749710), .ZN(n25801) );
  XNOR2_X1 U20726 ( .A(n24287), .B(n25794), .ZN(n25796) );
  NAND2_X1 U20727 ( .A1(n24322), .A2(net749822), .ZN(n26157) );
  NAND2_X1 U20728 ( .A1(net749312), .A2(net716215), .ZN(n25861) );
  NAND2_X1 U20729 ( .A1(n25789), .A2(n26027), .ZN(n26531) );
  NOR2_X1 U20730 ( .A1(net716237), .A2(\core_inst/EXMEM_NPC/DFF_12/N3 ), .ZN(
        n25470) );
  NOR2_X1 U20731 ( .A1(net749894), .A2(n25461), .ZN(n25460) );
  NAND2_X1 U20732 ( .A1(n26210), .A2(net713736), .ZN(n25459) );
  AND2_X1 U20733 ( .A1(\core_inst/MEM/MUX_LOAD/MUX_BIT_3/s_top ), .A2(n18200), 
        .ZN(\core_inst/MEMWB_DATAOUT/DFF_3/N3 ) );
  AND2_X1 U20734 ( .A1(\core_inst/MEM/MUX_LOAD/MUX_BIT_7/s_top ), .A2(n18200), 
        .ZN(\core_inst/MEMWB_DATAOUT/DFF_7/N3 ) );
  AND2_X1 U20735 ( .A1(\core_inst/MEM/MUX_LOAD/MUX_BIT_6/s_top ), .A2(n18200), 
        .ZN(\core_inst/MEMWB_DATAOUT/DFF_6/N3 ) );
  AND2_X1 U20736 ( .A1(\core_inst/MEM/MUX_LOAD/MUX_BIT_5/s_top ), .A2(n18200), 
        .ZN(\core_inst/MEMWB_DATAOUT/DFF_5/N3 ) );
  AND2_X1 U20737 ( .A1(\core_inst/MEM/MUX_LOAD/MUX_BIT_4/s_top ), .A2(n18200), 
        .ZN(\core_inst/MEMWB_DATAOUT/DFF_4/N3 ) );
  AND2_X1 U20738 ( .A1(\core_inst/MEM/MUX_LOAD/MUX_BIT_2/s_top ), .A2(n18200), 
        .ZN(\core_inst/MEMWB_DATAOUT/DFF_2/N3 ) );
  AND2_X1 U20739 ( .A1(\core_inst/MEM/MUX_LOAD/MUX_BIT_1/s_top ), .A2(n18200), 
        .ZN(\core_inst/MEMWB_DATAOUT/DFF_1/N3 ) );
  NOR2_X1 U20740 ( .A1(n26778), .A2(n20067), .ZN(n25666) );
  NOR2_X1 U20741 ( .A1(n26778), .A2(n20067), .ZN(n19351) );
  NAND2_X1 U20742 ( .A1(net755097), .A2(net742326), .ZN(n26018) );
  AOI22_X1 U20743 ( .A1(net713845), .A2(\core_inst/MEMWB_ALUOUT/DFF_16/N3 ), 
        .B1(net717789), .B2(n952), .ZN(n26048) );
  OAI22_X1 U20744 ( .A1(net717106), .A2(n1712), .B1(net714943), .B2(n25347), 
        .ZN(n25842) );
  OAI22_X1 U20745 ( .A1(net749972), .A2(n1748), .B1(net714943), .B2(n4416), 
        .ZN(n25829) );
  NAND3_X1 U20746 ( .A1(net726959), .A2(n25472), .A3(net726961), .ZN(n25372)
         );
  NOR2_X1 U20747 ( .A1(n25373), .A2(net715048), .ZN(n26256) );
  NOR2_X1 U20748 ( .A1(n26057), .A2(n25376), .ZN(n25497) );
  NOR2_X1 U20749 ( .A1(n25374), .A2(net714267), .ZN(n25375) );
  AOI21_X1 U20750 ( .B1(n26028), .B2(net714306), .A(n25375), .ZN(n25907) );
  OAI211_X1 U20751 ( .C1(net742157), .C2(n25381), .A(n25488), .B(n25489), .ZN(
        n25486) );
  NAND3_X1 U20752 ( .A1(n25381), .A2(net713683), .A3(n25798), .ZN(n25799) );
  NOR2_X1 U20753 ( .A1(net741958), .A2(n4406), .ZN(n25841) );
  NAND4_X1 U20754 ( .A1(net742042), .A2(n24264), .A3(net749334), .A4(n26097), 
        .ZN(n26104) );
  NAND3_X1 U20755 ( .A1(net749289), .A2(net755137), .A3(n25982), .ZN(n25978)
         );
  NAND2_X1 U20756 ( .A1(n25397), .A2(net742286), .ZN(n25427) );
  NOR2_X1 U20757 ( .A1(n25391), .A2(n22686), .ZN(n25399) );
  OAI22_X1 U20758 ( .A1(n1746), .A2(net715419), .B1(n4412), .B2(net717719), 
        .ZN(n25401) );
  NAND2_X1 U20759 ( .A1(n24569), .A2(n18052), .ZN(n25753) );
  NAND2_X1 U20760 ( .A1(n24295), .A2(n25344), .ZN(n26049) );
  NAND2_X1 U20761 ( .A1(n26147), .A2(n24572), .ZN(n26153) );
  OAI22_X1 U20762 ( .A1(net731327), .A2(net728314), .B1(net717075), .B2(
        net742259), .ZN(n25464) );
  OAI22_X1 U20763 ( .A1(net717875), .A2(n24357), .B1(net796212), .B2(net742324), .ZN(n25877) );
  AOI22_X1 U20764 ( .A1(n23022), .A2(net750032), .B1(n22948), .B2(net780543), 
        .ZN(n25808) );
  NAND2_X1 U20765 ( .A1(n24309), .A2(n24830), .ZN(n25422) );
  MUX2_X1 U20766 ( .A(n26171), .B(n26170), .S(net734022), .Z(net713762) );
  NOR2_X1 U20767 ( .A1(net714476), .A2(n24566), .ZN(n26059) );
  NOR2_X1 U20768 ( .A1(net742100), .A2(net754997), .ZN(n26731) );
  OAI22_X1 U20769 ( .A1(net742315), .A2(net762754), .B1(n24546), .B2(net713868), .ZN(n25951) );
  OAI22_X1 U20770 ( .A1(net742508), .A2(net717059), .B1(net717056), .B2(n25578), .ZN(n25463) );
  NOR2_X1 U20771 ( .A1(net742198), .A2(n23030), .ZN(n26739) );
  NAND2_X1 U20772 ( .A1(n25845), .A2(n26212), .ZN(n25936) );
  NAND3_X1 U20773 ( .A1(n25578), .A2(net742339), .A3(n22673), .ZN(n26044) );
  NAND2_X1 U20774 ( .A1(n24567), .A2(net755214), .ZN(n25781) );
  AOI22_X1 U20775 ( .A1(net717875), .A2(net765429), .B1(n22949), .B2(net714249), .ZN(n25433) );
  NAND2_X1 U20776 ( .A1(net718391), .A2(net765429), .ZN(n26045) );
  NAND2_X1 U20777 ( .A1(n24577), .A2(net750057), .ZN(n26024) );
  NAND2_X1 U20778 ( .A1(n25417), .A2(net713753), .ZN(n25856) );
  NAND2_X1 U20779 ( .A1(n25417), .A2(net749387), .ZN(n25761) );
  OAI21_X1 U20780 ( .B1(net713602), .B2(n22836), .A(net749465), .ZN(n25777) );
  MUX2_X1 U20781 ( .A(n25997), .B(n25419), .S(net717510), .Z(net714401) );
  OAI22_X1 U20782 ( .A1(net750278), .A2(net742087), .B1(net785220), .B2(
        net713773), .ZN(n25465) );
  NOR3_X1 U20783 ( .A1(n24310), .A2(net717875), .A3(net767203), .ZN(n25474) );
  OAI222_X1 U20784 ( .A1(n24310), .A2(net718391), .B1(net717055), .B2(n25586), 
        .C1(n24291), .C2(net742087), .ZN(n25954) );
  NAND2_X1 U20785 ( .A1(n22834), .A2(n25426), .ZN(n26066) );
  NAND3_X1 U20786 ( .A1(n24098), .A2(net713775), .A3(net755134), .ZN(n25476)
         );
  NAND3_X1 U20787 ( .A1(n25959), .A2(n25428), .A3(n24536), .ZN(net714261) );
  NAND2_X1 U20788 ( .A1(n24577), .A2(n26148), .ZN(n25434) );
  MUX2_X1 U20789 ( .A(net713728), .B(net713770), .S(n26223), .Z(n25436) );
  MUX2_X1 U20790 ( .A(net713726), .B(n25662), .S(n26223), .Z(n25435) );
  NAND3_X1 U20791 ( .A1(n25432), .A2(n25433), .A3(n25434), .ZN(n25431) );
  MUX2_X1 U20792 ( .A(n25435), .B(n25436), .S(n24311), .Z(n25430) );
  OAI211_X1 U20793 ( .C1(n25429), .C2(net739078), .A(n25430), .B(n25431), .ZN(
        net714241) );
  NAND2_X1 U20794 ( .A1(n25437), .A2(net742286), .ZN(n25934) );
  OAI22_X1 U20795 ( .A1(net755699), .A2(n24270), .B1(n24546), .B2(net742087), 
        .ZN(n25929) );
  OAI22_X1 U20796 ( .A1(net742483), .A2(n24546), .B1(n24270), .B2(n24269), 
        .ZN(n25911) );
  NAND2_X1 U20797 ( .A1(n25443), .A2(n24233), .ZN(n25790) );
  OAI22_X1 U20798 ( .A1(n24358), .A2(n24546), .B1(n24233), .B2(net742271), 
        .ZN(n25878) );
  NAND2_X1 U20799 ( .A1(n25450), .A2(n25451), .ZN(n25448) );
  AOI21_X1 U20800 ( .B1(n26023), .B2(net742339), .A(n24300), .ZN(n25450) );
  MUX2_X1 U20801 ( .A(net713892), .B(n26136), .S(n26210), .Z(n25461) );
  OAI22_X1 U20802 ( .A1(net713894), .A2(net714382), .B1(net713897), .B2(
        net714401), .ZN(n25456) );
  OAI222_X1 U20803 ( .A1(n26211), .A2(net713728), .B1(net713882), .B2(n26135), 
        .C1(net749977), .C2(net713977), .ZN(n25454) );
  OAI22_X1 U20804 ( .A1(net786856), .A2(net750287), .B1(n24560), .B2(net713810), .ZN(n25462) );
  MUX2_X1 U20805 ( .A(n25459), .B(n25460), .S(net755740), .Z(n25458) );
  NOR2_X1 U20806 ( .A1(n26581), .A2(net742182), .ZN(n26727) );
  NAND3_X1 U20807 ( .A1(n24203), .A2(net713775), .A3(net750090), .ZN(n25477)
         );
  NAND3_X1 U20808 ( .A1(n24355), .A2(net713775), .A3(net714194), .ZN(n25484)
         );
  NAND3_X1 U20809 ( .A1(net713748), .A2(net713775), .A3(n26064), .ZN(n25483)
         );
  NAND3_X1 U20810 ( .A1(net712466), .A2(net713775), .A3(net713707), .ZN(n25482) );
  NAND3_X1 U20811 ( .A1(net712468), .A2(net713775), .A3(n26071), .ZN(n25481)
         );
  NAND3_X1 U20812 ( .A1(n24340), .A2(net713775), .A3(n24359), .ZN(n25489) );
  NAND3_X1 U20813 ( .A1(n24550), .A2(net713775), .A3(net780543), .ZN(n25488)
         );
  NAND3_X1 U20814 ( .A1(n24556), .A2(net713775), .A3(net749732), .ZN(n25493)
         );
  MUX2_X1 U20815 ( .A(n25494), .B(n25495), .S(net742157), .Z(n25492) );
  NAND2_X1 U20816 ( .A1(n25501), .A2(n24548), .ZN(n25499) );
  NAND3_X1 U20817 ( .A1(n26054), .A2(n26056), .A3(net739078), .ZN(n25498) );
  NOR3_X1 U20818 ( .A1(net767203), .A2(n24577), .A3(net717074), .ZN(n25479) );
  NOR3_X1 U20819 ( .A1(n26063), .A2(net762661), .A3(net767203), .ZN(n25487) );
  NAND3_X1 U20820 ( .A1(n25498), .A2(n25499), .A3(n25500), .ZN(n25496) );
  AOI211_X1 U20821 ( .C1(n25473), .C2(n24566), .A(n25474), .B(n25475), .ZN(
        net714175) );
  NOR4_X1 U20822 ( .A1(n25485), .A2(n25486), .A3(n25316), .A4(n25487), .ZN(
        net714173) );
  NOR2_X1 U20823 ( .A1(n25496), .A2(n25497), .ZN(net714172) );
  XNOR2_X1 U20824 ( .A(n25995), .B(net716215), .ZN(n25835) );
  NAND2_X1 U20825 ( .A1(n25835), .A2(net714494), .ZN(n25992) );
  NAND3_X1 U20826 ( .A1(n25752), .A2(net786837), .A3(net725586), .ZN(n25508)
         );
  NAND3_X1 U20827 ( .A1(n25758), .A2(n26185), .A3(n25757), .ZN(n25510) );
  OAI21_X1 U20828 ( .B1(net716333), .B2(n25536), .A(n25537), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_26/N3 ) );
  OAI21_X1 U20829 ( .B1(net796193), .B2(n25544), .A(n25545), .ZN(
        \core_inst/IDEX_RF_IN1/DFF_14/N3 ) );
  OAI21_X1 U20830 ( .B1(net716313), .B2(n25557), .A(n25558), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_21/N3 ) );
  OAI21_X1 U20831 ( .B1(net796133), .B2(n25549), .A(n25550), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_29/N3 ) );
  OAI21_X1 U20832 ( .B1(net796133), .B2(n25565), .A(n25566), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_4/N3 ) );
  OAI21_X1 U20833 ( .B1(net716369), .B2(n25569), .A(n25570), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_18/N3 ) );
  NAND3_X1 U20834 ( .A1(net716263), .A2(net717050), .A3(n26652), .ZN(n25558)
         );
  NAND3_X1 U20835 ( .A1(net716265), .A2(net717050), .A3(n26718), .ZN(n25566)
         );
  NAND3_X1 U20836 ( .A1(net742368), .A2(net717049), .A3(n26706), .ZN(n25570)
         );
  NOR2_X1 U20837 ( .A1(net716333), .A2(n5596), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_29/N3 ) );
  NOR2_X1 U20838 ( .A1(net812952), .A2(n371), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_25/N3 ) );
  NOR2_X1 U20839 ( .A1(net796193), .A2(n562), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_27/N3 ) );
  OAI22_X1 U20840 ( .A1(net713773), .A2(n24559), .B1(n24233), .B2(n25578), 
        .ZN(n25950) );
  OAI22_X1 U20841 ( .A1(net731327), .A2(net796212), .B1(net755757), .B2(
        net718355), .ZN(n26121) );
  AND2_X1 U20842 ( .A1(\core_inst/MEM/MUX_LOAD/MUX_BIT_0/s_top ), .A2(n18200), 
        .ZN(\core_inst/MEMWB_DATAOUT/DFF_0/N3 ) );
  OAI21_X1 U20843 ( .B1(n25800), .B2(net713683), .A(n25799), .ZN(n25802) );
  NAND2_X1 U20844 ( .A1(net712466), .A2(net713683), .ZN(n25806) );
  AOI21_X1 U20845 ( .B1(n25932), .B2(n25931), .A(net713751), .ZN(n25933) );
  NAND2_X1 U20846 ( .A1(n24547), .A2(n25994), .ZN(n26192) );
  NAND2_X1 U20847 ( .A1(n24577), .A2(n24280), .ZN(n26191) );
  NOR2_X1 U20848 ( .A1(net716311), .A2(net762759), .ZN(
        \core_inst/EXMEM_IR/DFF_20/N3 ) );
  NOR2_X1 U20849 ( .A1(net796193), .A2(n24581), .ZN(
        \core_inst/IDEX_IR/DFF_27/N3 ) );
  AOI21_X1 U20850 ( .B1(n6402), .B2(net712838), .A(n26457), .ZN(n26458) );
  NAND2_X1 U20851 ( .A1(n24561), .A2(net749710), .ZN(n25817) );
  NOR2_X1 U20852 ( .A1(net765727), .A2(n24534), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_2/N3 ) );
  NOR2_X1 U20853 ( .A1(n26727), .A2(net796232), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_20/N3 ) );
  NOR2_X1 U20854 ( .A1(net812279), .A2(n17689), .ZN(
        \core_inst/IDEX_NPC/DFF_25/N3 ) );
  NOR2_X1 U20855 ( .A1(net804592), .A2(n6555), .ZN(
        \core_inst/IDEX_NPC/DFF_9/N3 ) );
  NOR2_X1 U20856 ( .A1(net785270), .A2(n26730), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_13/N3 ) );
  NOR2_X1 U20857 ( .A1(net765319), .A2(n26729), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_15/N3 ) );
  NOR2_X1 U20858 ( .A1(net812958), .A2(n26728), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_16/N3 ) );
  NOR2_X1 U20859 ( .A1(net804592), .A2(net712390), .ZN(
        \core_inst/EXMEM_IR/DFF_29/N3 ) );
  NOR2_X1 U20860 ( .A1(net796193), .A2(n24785), .ZN(
        \core_inst/IDEX_IMM_IN/DFF_4/N3 ) );
  NOR2_X1 U20861 ( .A1(net716353), .A2(n1539), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_0/N3 ) );
  NOR2_X1 U20862 ( .A1(net796114), .A2(n6475), .ZN(
        \core_inst/IDEX_NPC/DFF_2/N3 ) );
  NOR2_X1 U20863 ( .A1(net796193), .A2(n26731), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_9/N3 ) );
  NOR2_X1 U20864 ( .A1(net716313), .A2(n5602), .ZN(
        \core_inst/EXMEM_DATAIN/DFF_28/N3 ) );
  NOR2_X1 U20865 ( .A1(net796143), .A2(n1222), .ZN(
        \core_inst/IDEX_NPC/DFF_10/N3 ) );
  NOR2_X1 U20866 ( .A1(net716311), .A2(n26732), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_18/N3 ) );
  NOR2_X1 U20867 ( .A1(net716311), .A2(n26734), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_26/N3 ) );
  NOR2_X1 U20868 ( .A1(net716313), .A2(n26736), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_22/N3 ) );
  NOR2_X1 U20869 ( .A1(net716353), .A2(n26735), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_30/N3 ) );
  OAI21_X1 U20870 ( .B1(n26731), .B2(net716267), .A(n26707), .ZN(n16391) );
  OAI21_X1 U20871 ( .B1(n26734), .B2(net716263), .A(n26711), .ZN(n26783) );
  OAI21_X1 U20872 ( .B1(n26730), .B2(net765341), .A(n26713), .ZN(n26784) );
  NOR2_X1 U20873 ( .A1(n25881), .A2(n25880), .ZN(n25882) );
  NOR2_X1 U20874 ( .A1(net716333), .A2(net718087), .ZN(
        \core_inst/EXMEM_IR/DFF_16/N3 ) );
  AOI21_X1 U20875 ( .B1(n6746), .B2(n1498), .A(n26604), .ZN(n26744) );
  AOI21_X1 U20876 ( .B1(n5171), .B2(n26558), .A(net785319), .ZN(n26559) );
  AOI21_X1 U20877 ( .B1(n6511), .B2(n26578), .A(net712922), .ZN(n26534) );
  AOI21_X1 U20878 ( .B1(n6516), .B2(net712490), .A(n26579), .ZN(n26530) );
  NAND4_X1 U20879 ( .A1(n22869), .A2(n24092), .A3(n26079), .A4(net749308), 
        .ZN(n26083) );
  NOR2_X1 U20880 ( .A1(net716313), .A2(net749817), .ZN(
        \core_inst/EXMEM_IR/DFF_17/N3 ) );
  AOI22_X1 U20881 ( .A1(n26164), .A2(n26167), .B1(net718391), .B2(net713748), 
        .ZN(net713760) );
  AOI22_X1 U20882 ( .A1(net712468), .A2(net714194), .B1(net712467), .B2(
        net750090), .ZN(n25809) );
  NAND4_X1 U20883 ( .A1(n24533), .A2(n26007), .A3(n26011), .A4(n26015), .ZN(
        net714463) );
  AOI22_X1 U20884 ( .A1(n26137), .A2(net713779), .B1(net713870), .B2(net713874), .ZN(n26016) );
  NAND2_X1 U20885 ( .A1(n24090), .A2(n24282), .ZN(n26563) );
  NAND2_X1 U20886 ( .A1(net755240), .A2(n25991), .ZN(n26230) );
  NAND2_X1 U20887 ( .A1(net713985), .A2(n26051), .ZN(n26053) );
  NOR2_X1 U20888 ( .A1(net716311), .A2(n24583), .ZN(
        \core_inst/IDEX_IR/DFF_29/N3 ) );
  XNOR2_X1 U20889 ( .A(n25793), .B(net713683), .ZN(n25794) );
  NAND2_X1 U20890 ( .A1(net748269), .A2(net739078), .ZN(n26218) );
  OAI22_X1 U20891 ( .A1(net749260), .A2(net762754), .B1(net717074), .B2(
        net748269), .ZN(n25797) );
  OAI22_X1 U20892 ( .A1(net742259), .A2(net762754), .B1(net717055), .B2(
        net755699), .ZN(n26122) );
  NOR2_X1 U20893 ( .A1(net716377), .A2(n26724), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_1/N3 ) );
  OAI21_X1 U20894 ( .B1(n26724), .B2(net716257), .A(net712391), .ZN(
        \core_inst/IF_stage/PROGRAM_COUNTER/DFF_1/N3 ) );
  OAI222_X1 U20895 ( .A1(n24342), .A2(net714182), .B1(net713154), .B2(n25864), 
        .C1(net714267), .C2(n26173), .ZN(n25870) );
  NAND2_X1 U20896 ( .A1(n24532), .A2(n24540), .ZN(n26092) );
  NOR2_X1 U20897 ( .A1(n25937), .A2(n25938), .ZN(n26131) );
  NOR2_X1 U20898 ( .A1(net762754), .A2(net742087), .ZN(n26004) );
  NOR2_X1 U20899 ( .A1(net785239), .A2(n24126), .ZN(
        \core_inst/EXMEM_ALU_OUT/DFF_6/N3 ) );
  NOR2_X1 U20900 ( .A1(n25957), .A2(n25958), .ZN(n25965) );
  OAI21_X1 U20901 ( .B1(net716313), .B2(n26660), .A(n26659), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_24/N3 ) );
  OAI21_X1 U20902 ( .B1(net812941), .B2(n26281), .A(n26280), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_23/N3 ) );
  NOR2_X1 U20903 ( .A1(n25938), .A2(net755139), .ZN(n25823) );
  AOI22_X1 U20904 ( .A1(n26039), .A2(net767208), .B1(n25594), .B2(net714275), 
        .ZN(n25819) );
  NAND2_X1 U20905 ( .A1(n25594), .A2(net714306), .ZN(n25968) );
  OAI21_X1 U20906 ( .B1(net796136), .B2(n26438), .A(n26437), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_27/N3 ) );
  OAI22_X1 U20907 ( .A1(net749343), .A2(net762754), .B1(net750287), .B2(
        net718391), .ZN(n25926) );
  OAI22_X1 U20908 ( .A1(net749454), .A2(net750287), .B1(n26063), .B2(net713810), .ZN(n25953) );
  NAND2_X1 U20909 ( .A1(n24191), .A2(net749454), .ZN(n25943) );
  AOI21_X1 U20910 ( .B1(n25956), .B2(n25955), .A(net713751), .ZN(n25957) );
  NOR2_X1 U20911 ( .A1(net712931), .A2(n26529), .ZN(n26729) );
  OAI22_X1 U20912 ( .A1(net749306), .A2(n24357), .B1(net796212), .B2(net749812), .ZN(n25910) );
  NAND2_X1 U20913 ( .A1(net749967), .A2(n25909), .ZN(n26156) );
  NAND2_X1 U20914 ( .A1(net750025), .A2(net742507), .ZN(n25857) );
  NAND2_X1 U20915 ( .A1(n25998), .A2(net749910), .ZN(n26154) );
  NAND2_X1 U20916 ( .A1(n25987), .A2(net749910), .ZN(n25783) );
  NAND2_X1 U20917 ( .A1(net762660), .A2(net717510), .ZN(n26217) );
  NAND2_X1 U20918 ( .A1(n24033), .A2(n23974), .ZN(n26196) );
  OAI22_X1 U20919 ( .A1(net750238), .A2(net728314), .B1(net796212), .B2(
        net750019), .ZN(n25949) );
  AOI22_X1 U20920 ( .A1(net718380), .A2(n24293), .B1(net750019), .B2(n24201), 
        .ZN(n26202) );
  NOR2_X1 U20921 ( .A1(n24177), .A2(net742242), .ZN(n26054) );
  NAND2_X1 U20922 ( .A1(net713754), .A2(net742243), .ZN(n26219) );
  NAND2_X1 U20923 ( .A1(net713677), .A2(net762625), .ZN(n25787) );
  NAND2_X1 U20924 ( .A1(net749612), .A2(n24192), .ZN(n26036) );
  OAI21_X1 U20925 ( .B1(n24534), .B2(net716267), .A(n26719), .ZN(
        \core_inst/IF_stage/PROGRAM_COUNTER/DFF_2/N3 ) );
  OAI21_X1 U20926 ( .B1(n26738), .B2(net742648), .A(n26716), .ZN(
        \core_inst/IF_stage/PROGRAM_COUNTER/DFF_11/N3 ) );
  OAI21_X1 U20927 ( .B1(n26695), .B2(n26694), .A(net716257), .ZN(n26696) );
  OAI22_X1 U20928 ( .A1(net717875), .A2(net750287), .B1(n26063), .B2(n24358), 
        .ZN(n25914) );
  NOR2_X1 U20929 ( .A1(net750228), .A2(net762597), .ZN(n26182) );
  OAI21_X1 U20930 ( .B1(n26322), .B2(n26321), .A(net741999), .ZN(n26323) );
  OAI21_X1 U20931 ( .B1(n26301), .B2(n26300), .A(net716247), .ZN(n26302) );
  OAI21_X1 U20932 ( .B1(n26391), .B2(n26390), .A(net742648), .ZN(n26392) );
  OAI21_X1 U20933 ( .B1(n26402), .B2(n26401), .A(net785255), .ZN(n26403) );
  OAI21_X1 U20934 ( .B1(n26311), .B2(n26310), .A(net716247), .ZN(n26312) );
  OAI21_X1 U20935 ( .B1(net796193), .B2(n26351), .A(n26350), .ZN(
        \core_inst/IDEX_RF_IN2/DFF_17/N3 ) );
  AOI211_X1 U20936 ( .C1(n25902), .C2(n24566), .A(n25901), .B(n25316), .ZN(
        n25908) );
  NAND2_X1 U20937 ( .A1(n25989), .A2(n24566), .ZN(n25946) );
  NAND2_X1 U20938 ( .A1(net716249), .A2(s_IFID_IR[19]), .ZN(n26577) );
  OAI21_X1 U20939 ( .B1(n26492), .B2(n26491), .A(net741999), .ZN(n26493) );
  OAI21_X1 U20940 ( .B1(n26650), .B2(n26649), .A(net716257), .ZN(n26651) );
  OAI21_X1 U20941 ( .B1(n26518), .B2(net712945), .A(net741999), .ZN(n26519) );
  OAI21_X1 U20942 ( .B1(n26480), .B2(n26479), .A(net716261), .ZN(n26481) );
  OAI21_X1 U20943 ( .B1(n26419), .B2(n26418), .A(net716261), .ZN(n26420) );
  OAI21_X1 U20944 ( .B1(n26469), .B2(n26468), .A(net760161), .ZN(n26470) );
  OAI22_X1 U20945 ( .A1(n24566), .A2(n26064), .B1(n24554), .B2(net717570), 
        .ZN(n25778) );
  NOR2_X1 U20946 ( .A1(net767341), .A2(n25357), .ZN(n25830) );
  NAND2_X1 U20947 ( .A1(net713677), .A2(n24206), .ZN(n26216) );
  NOR3_X1 U20948 ( .A1(n25954), .A2(n25953), .A3(n25952), .ZN(n25955) );
  NAND2_X1 U20949 ( .A1(net755238), .A2(net714249), .ZN(n26025) );
  NAND2_X1 U20950 ( .A1(net713773), .A2(net714249), .ZN(n26043) );
  OAI22_X1 U20951 ( .A1(net742507), .A2(n25599), .B1(net713907), .B2(net713905), .ZN(n25952) );
  OAI22_X1 U20952 ( .A1(n25586), .A2(n24357), .B1(net796212), .B2(net750238), 
        .ZN(n25928) );
  NAND2_X1 U20953 ( .A1(n25586), .A2(n24198), .ZN(n26206) );
  NAND2_X1 U20954 ( .A1(net749898), .A2(net713810), .ZN(n26155) );
  NAND2_X1 U20955 ( .A1(net749489), .A2(net749387), .ZN(n25858) );
  NOR2_X1 U20956 ( .A1(net718351), .A2(n953), .ZN(n25849) );
  NAND3_X1 U20957 ( .A1(n25779), .A2(net717510), .A3(n25393), .ZN(net712893)
         );
  MUX2_X1 U20958 ( .A(net767234), .B(net713736), .S(net713554), .Z(n26408) );
  MUX2_X1 U20959 ( .A(net767234), .B(net713736), .S(net742092), .Z(n25800) );
  MUX2_X1 U20960 ( .A(net713726), .B(net713738), .S(net742092), .Z(n25798) );
  NAND3_X1 U20961 ( .A1(n25803), .A2(n25802), .A3(n25801), .ZN(n25804) );
  MUX2_X1 U20962 ( .A(net713726), .B(n25662), .S(n25816), .Z(n25810) );
  MUX2_X1 U20963 ( .A(n25812), .B(n25811), .S(n26064), .Z(n25813) );
  XOR2_X1 U20964 ( .A(n24358), .B(n24564), .Z(n25863) );
  XOR2_X1 U20965 ( .A(n25863), .B(n25862), .Z(n25864) );
  MUX2_X1 U20966 ( .A(net713726), .B(net713738), .S(n25579), .Z(n25865) );
  MUX2_X1 U20967 ( .A(net767234), .B(net713736), .S(n25579), .Z(n25866) );
  MUX2_X1 U20968 ( .A(n25867), .B(n25866), .S(n24358), .Z(n25868) );
  MUX2_X1 U20969 ( .A(net713726), .B(net713728), .S(net713753), .Z(n25889) );
  MUX2_X1 U20970 ( .A(n25662), .B(net713770), .S(net713753), .Z(n25888) );
  MUX2_X1 U20971 ( .A(n25889), .B(n25888), .S(n26194), .Z(n25890) );
  MUX2_X1 U20972 ( .A(net713728), .B(net713726), .S(n24548), .Z(n25905) );
  MUX2_X1 U20973 ( .A(net713770), .B(net713738), .S(n24548), .Z(n25904) );
  MUX2_X1 U20974 ( .A(n25905), .B(n25904), .S(n23966), .Z(n25906) );
  NAND3_X1 U20975 ( .A1(n25908), .A2(n25907), .A3(n25906), .ZN(n25919) );
  MUX2_X1 U20976 ( .A(n26047), .B(n25947), .S(net718367), .Z(n25958) );
  MUX2_X1 U20977 ( .A(net767234), .B(net713736), .S(n23974), .Z(n25960) );
  MUX2_X1 U20978 ( .A(n25961), .B(n25960), .S(n24341), .Z(n25962) );
  MUX2_X1 U20979 ( .A(net713728), .B(net713726), .S(net713707), .Z(n25967) );
  MUX2_X1 U20980 ( .A(net717087), .B(net713738), .S(net713707), .Z(n25966) );
  MUX2_X1 U20981 ( .A(n25967), .B(n25966), .S(n24285), .Z(n25969) );
  NAND3_X1 U20982 ( .A1(n26072), .A2(net714603), .A3(n25976), .ZN(n25977) );
  MUX2_X1 U20983 ( .A(n25988), .B(n25987), .S(net742339), .Z(n26000) );
  MUX2_X1 U20984 ( .A(net713892), .B(n26136), .S(n26228), .Z(n26003) );
  MUX2_X1 U20985 ( .A(net767234), .B(net713736), .S(n26228), .Z(n26002) );
  MUX2_X1 U20986 ( .A(n26003), .B(n26002), .S(net786856), .Z(n26010) );
  NAND3_X1 U20987 ( .A1(n26016), .A2(n26017), .A3(n26015), .ZN(net714466) );
  NAND3_X1 U20988 ( .A1(n26095), .A2(n26094), .A3(n26093), .ZN(net714033) );
  NAND3_X1 U20989 ( .A1(n26117), .A2(n26116), .A3(n26115), .ZN(net714034) );
  NAND3_X1 U20990 ( .A1(n26125), .A2(n26124), .A3(n26123), .ZN(n26126) );
  MUX2_X1 U20991 ( .A(net713892), .B(n26136), .S(net762674), .Z(n26133) );
  MUX2_X1 U20992 ( .A(n26146), .B(n26145), .S(net750176), .Z(n26147) );
  NAND3_X1 U20993 ( .A1(net742157), .A2(n26148), .A3(net749534), .ZN(n26151)
         );
  NAND3_X1 U20994 ( .A1(n26158), .A2(net713785), .A3(n26157), .ZN(n26159) );
  MUX2_X1 U20995 ( .A(net713738), .B(net713726), .S(n26168), .Z(n26169) );
  NAND3_X1 U20996 ( .A1(n26189), .A2(n26188), .A3(net750090), .ZN(n26237) );
  NAND3_X1 U20997 ( .A1(net716247), .A2(net717050), .A3(n26478), .ZN(n26280)
         );
  NAND3_X1 U20998 ( .A1(n26287), .A2(n26286), .A3(n26285), .ZN(n26288) );
  NAND3_X1 U20999 ( .A1(n19145), .A2(n19146), .A3(n26291), .ZN(n26293) );
  NAND3_X1 U21000 ( .A1(n19161), .A2(n19160), .A3(n19159), .ZN(n26292) );
  NAND3_X1 U21001 ( .A1(n26294), .A2(n19165), .A3(n19158), .ZN(n26296) );
  NAND3_X1 U21002 ( .A1(n19520), .A2(n19521), .A3(n26303), .ZN(n26308) );
  NAND3_X1 U21003 ( .A1(n19537), .A2(n19531), .A3(n19536), .ZN(n26306) );
  NAND3_X1 U21004 ( .A1(n19534), .A2(n19533), .A3(n19532), .ZN(n26305) );
  NAND3_X1 U21005 ( .A1(n19232), .A2(n19233), .A3(n26313), .ZN(n26315) );
  NAND3_X1 U21006 ( .A1(n19269), .A2(n19268), .A3(n19267), .ZN(n26314) );
  NAND3_X1 U21007 ( .A1(n26316), .A2(n19275), .A3(n19266), .ZN(n26318) );
  NAND3_X1 U21008 ( .A1(n19873), .A2(n19874), .A3(n26324), .ZN(n26326) );
  NAND3_X1 U21009 ( .A1(n19631), .A2(n19632), .A3(n26329), .ZN(n26332) );
  NAND3_X1 U21010 ( .A1(n19609), .A2(n19610), .A3(n26352), .ZN(n26357) );
  NAND3_X1 U21011 ( .A1(n19625), .A2(n19619), .A3(n19624), .ZN(n26355) );
  NAND3_X1 U21012 ( .A1(n19622), .A2(n19621), .A3(n19620), .ZN(n26354) );
  NAND3_X1 U21013 ( .A1(n19510), .A2(n19509), .A3(n19508), .ZN(n26360) );
  NAND3_X1 U21014 ( .A1(n19173), .A2(n19174), .A3(n26374), .ZN(n26376) );
  NAND3_X1 U21015 ( .A1(n19189), .A2(n19188), .A3(n19187), .ZN(n26375) );
  NAND3_X1 U21016 ( .A1(n26377), .A2(n19193), .A3(n19186), .ZN(n26379) );
  NAND3_X1 U21017 ( .A1(n19587), .A2(n19588), .A3(n26383), .ZN(n26388) );
  NAND3_X1 U21018 ( .A1(n19603), .A2(n19597), .A3(n19602), .ZN(n26386) );
  NAND3_X1 U21019 ( .A1(n19600), .A2(n19599), .A3(n19598), .ZN(n26385) );
  NAND3_X1 U21020 ( .A1(n19851), .A2(n19852), .A3(n26393), .ZN(n26398) );
  NAND3_X1 U21021 ( .A1(n19867), .A2(n19861), .A3(n19866), .ZN(n26396) );
  NAND3_X1 U21022 ( .A1(n19864), .A2(n19863), .A3(n19862), .ZN(n26395) );
  NAND3_X1 U21023 ( .A1(n19675), .A2(n19676), .A3(n26411), .ZN(n26416) );
  NAND3_X1 U21024 ( .A1(n19691), .A2(n19685), .A3(n19690), .ZN(n26414) );
  NAND3_X1 U21025 ( .A1(n19688), .A2(n19687), .A3(n19686), .ZN(n26413) );
  NAND3_X1 U21026 ( .A1(n19807), .A2(n19808), .A3(n26421), .ZN(n26426) );
  NAND3_X1 U21027 ( .A1(n19823), .A2(n19817), .A3(n19822), .ZN(n26424) );
  NAND3_X1 U21028 ( .A1(n19820), .A2(n19819), .A3(n19818), .ZN(n26423) );
  NAND3_X1 U21029 ( .A1(net742368), .A2(net712397), .A3(n26436), .ZN(n26437)
         );
  NAND3_X1 U21030 ( .A1(n20054), .A2(n20055), .A3(n26439), .ZN(n26446) );
  NAND3_X1 U21031 ( .A1(n20088), .A2(n20087), .A3(n20086), .ZN(n26444) );
  NAND3_X1 U21032 ( .A1(n19719), .A2(n19720), .A3(n26449), .ZN(n26454) );
  NAND3_X1 U21033 ( .A1(n19735), .A2(n19729), .A3(n19734), .ZN(n26452) );
  NAND3_X1 U21034 ( .A1(n19732), .A2(n19731), .A3(n19730), .ZN(n26451) );
  NAND3_X1 U21035 ( .A1(n19653), .A2(n19654), .A3(n26460), .ZN(n26465) );
  NAND3_X1 U21036 ( .A1(n19669), .A2(n19663), .A3(n19668), .ZN(n26463) );
  NAND3_X1 U21037 ( .A1(n19666), .A2(n19665), .A3(n19664), .ZN(n26462) );
  NAND3_X1 U21038 ( .A1(n19697), .A2(n19698), .A3(n26471), .ZN(n26476) );
  NAND3_X1 U21039 ( .A1(n19713), .A2(n19707), .A3(n19712), .ZN(n26474) );
  NAND3_X1 U21040 ( .A1(n19710), .A2(n19709), .A3(n19708), .ZN(n26473) );
  NAND3_X1 U21041 ( .A1(n19201), .A2(n19202), .A3(n26482), .ZN(n26484) );
  NAND3_X1 U21042 ( .A1(n19217), .A2(n19216), .A3(n19215), .ZN(n26483) );
  NAND3_X1 U21043 ( .A1(n26485), .A2(n19221), .A3(n19214), .ZN(n26487) );
  NAND3_X1 U21044 ( .A1(n19779), .A2(n19773), .A3(n19778), .ZN(n26514) );
  NAND3_X1 U21045 ( .A1(n19776), .A2(n19775), .A3(n19774), .ZN(n26513) );
  NAND3_X1 U21046 ( .A1(n19565), .A2(n19566), .A3(n26583), .ZN(n26588) );
  NAND3_X1 U21047 ( .A1(n19581), .A2(n19575), .A3(n19580), .ZN(n26586) );
  NAND3_X1 U21048 ( .A1(n19578), .A2(n19577), .A3(n19576), .ZN(n26585) );
  NAND3_X1 U21049 ( .A1(n26598), .A2(n26597), .A3(n26596), .ZN(n26599) );
  NAND3_X1 U21050 ( .A1(n20013), .A2(n20012), .A3(n20011), .ZN(n26627) );
  NAND3_X1 U21051 ( .A1(n19829), .A2(n19830), .A3(n26632), .ZN(n26636) );
  NAND3_X1 U21052 ( .A1(n19845), .A2(n19839), .A3(n19844), .ZN(n26634) );
  NAND3_X1 U21053 ( .A1(n19034), .A2(n19035), .A3(n26640), .ZN(n26642) );
  NAND3_X1 U21054 ( .A1(n19050), .A2(n19049), .A3(n19048), .ZN(n26641) );
  NAND3_X1 U21055 ( .A1(n26643), .A2(n19054), .A3(n19047), .ZN(n26645) );
  NAND3_X1 U21056 ( .A1(net716247), .A2(net717049), .A3(n26658), .ZN(n26659)
         );
  NAND3_X1 U21057 ( .A1(n18324), .A2(n18323), .A3(n18322), .ZN(n26682) );
  NAND3_X1 U21058 ( .A1(n19117), .A2(n19118), .A3(n26686), .ZN(n26688) );
  NAND3_X1 U21059 ( .A1(n19133), .A2(n19132), .A3(n19131), .ZN(n26687) );
  NAND3_X1 U21060 ( .A1(n26689), .A2(n19137), .A3(n19130), .ZN(n26691) );
  NAND3_X1 U21061 ( .A1(n26697), .A2(n19082), .A3(n19075), .ZN(n26699) );
endmodule

