library ieee;
use ieee.std_logic_1164.all;
use work.CU_pkg.all;

entity cu_core is
    generic(
        CU_IR_NBIT  :   positive    :=  32);
    port(
        CU_instruction_register :   in  std_logic_vector(CU_IR_NBIT-1 downto 0);
        CU_decode_ext_op        :   out std_logic_vector(1 downto 0);
        CU_decode_dest_sel      :   out std_logic;
        CU_execute_branch_type  :   out std_logic;
        CU_execute_alu_op       :   out std_logic_vector(5 downto 0);
        CU_execute_top_mux      :   out std_logic;
        CU_execute_bottom_mux   :   out std_logic;
        CU_execute_is_branch    :   out std_logic;
        CU_memory_r_not_w       :   out std_logic;
        CU_memory_signed_load   :   out std_logic;
        CU_memory_load_type     :   out std_logic_vector(1 downto 0);
        CU_writeback_write_en   :   out std_logic;
        CU_writeback_mux        :   out std_logic);
end entity;

architecture bhv of cu_core is

    signal s_cu_opcode(CU_OPCODE_NBIT-1 downto 0);
    signal s_cu_func(CU_FUNC_NBIT-1 downto 0);

begin

    s_cu_opcode <=  CU_instruction_register(CU_IR_NBIT-1 downto CU_IR_NBIT-CU_OPCODE_NBIT);
    s_cu_func   <=  CU_instruction_register(CU_FUNC_NBIT-1 downto 0);

    MAIN : process(CU_instruction_register)
    begin
        case(s_cu_opcode) is
            when CU_ALU_OPCODE =>
                case(s_cu_func) is
                    when sll        =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when srl        =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when sra        =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when add        =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when addu       =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when sub        =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when subu       =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when and        =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when or         =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when xor        =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when seq        =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when sne        =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when slt        =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when sgt        =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when sle        =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when sge        =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when sltu       =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when sgtu       =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when sleu       =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when sgeu       =>
                        CU_decode_signed_ext    <=
                        CU_execute_alu_op       <=
                        CU_execute_top_mux      <=
                        CU_execute_bottom_mux   <=
                        CU_memory_r_not_w       <=
                        CU_memory_signed_load   <=
                        CU_memory_load_type     <=
                        CU_writeback_write_en   <=
                        CU_writeback_mux        <=
                    when others     =>
                end case;
            when j      =>
                CU_decode_ext_op        <=  "01",       --  extend as 23 bits unsigned immediate
                CU_decode_dest_sel      <=  "00",       --  don't care
                CU_decode_read1_en      <=  '0',        --  don't read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '1',        --  j is always taken
                CU_execute_alu_op       <=  "010000"    --  add immediate target to 0
                CU_execute_top_mux      <=  '1',        --  read all zero from RF_in1
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '1',        --  is branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '0',        --  don't write anything
                CU_writeback_mux        <=  "00",       --  don't care
            when jal    =>
                CU_decode_ext_op        <=  "01",       --  extend as 23 bits unsigned immedaite
                CU_decode_dest_sel      <=  "11",       --  force register 31 as destination
                CU_decode_read1_en      <=  '0',        --  don't read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '1',        --  j is always taken
                CU_execute_alu_op       <=  "010000"    --  add immediate target to 0
                CU_execute_top_mux      <=  '1',        --  read all zero from RF_in1
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '1',        --  is branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write npc to register 31
                CU_writeback_mux        <=  "10"        --  write NPC
            when beqz   =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immedaite
                CU_decode_dest_sel      <=  "00",       --  don't care
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '1',        --  branch equal zero
                CU_execute_alu_op       <=  "010000"    --  add
                CU_execute_top_mux      <=  '0',        --  take NPC
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '1',        --  is branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '0',        --  don't write anything
                CU_writeback_mux        <=  "00"        --  don't write anything
            when bnez   =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immedaite
                CU_decode_dest_sel      <=  "00",       --  don't care
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  branch not equal zero
                CU_execute_alu_op       <=  "010000"    --  add
                CU_execute_top_mux      <=  '0',        --  take NPC
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '1',        --  is branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '0',        --  don't write anything
                CU_writeback_mux        <=  "00"        --  don't write anything
            when addi   =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immedaite
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '1',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "010000"    --  add
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "01"        --  write data from ALU
            when addui  =>
                CU_decode_ext_op        <=  "00",       --  extend as 16 bits unsigned immedaite
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '1',        --  read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "010000"    --  add
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "01"        --  write data from ALU
            when subi   =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immedaite
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '1',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "011000"    --  sub
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "01"        --  write data from ALU
            when subui  =>
                CU_decode_ext_op        <=  "00",       --  extend as 16 bits unsigned immedaite
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '1',        --  read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "011000"    --  sub
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "01"        --  write data from ALU
            when andi   =>
                CU_decode_ext_op        <=  "00",       --  extend as 16 bits unsigned immedaite
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '1',        --  read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "111000"    --  and
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "01"        --  write data from ALU
            when ori    =>
                CU_decode_ext_op        <=  "00",       --  extend as 16 bits unsigned immedaite
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '1',        --  read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "111110"    --  or
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "01"        --  write data from ALU
            when xori   =>
                CU_decode_ext_op        <=  "00",       --  extend as 16 bits unsigned immedaite
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '1',        --  read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "110110"    --  xor
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "01"        --  write data from ALU
            when lhi    =>  --  still to do
            when jr     =>
                CU_decode_ext_op        <=  "00",       --  don't care
                CU_decode_dest_sel      <=  "00",       --  don't care
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '1',        --  absolute branch
                CU_execute_alu_op       <=  "010000"    --  add
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  don't care
                CU_execute_is_branch    <=  '1',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '0',        --  write to rf
                CU_writeback_mux        <=  "00"        --  don't care
            when jalr   =>
                CU_decode_ext_op        <=  "00",       --  don't care
                CU_decode_dest_sel      <=  "11",       --  force register 31 as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '1',        --  j is always taken
                CU_execute_alu_op       <=  "010000"    --  add immediate target to 0
                CU_execute_top_mux      <=  '1',        --  read rs
                CU_execute_bottom_mux   <=  '1',        --  read all zero from RF_in2
                CU_execute_is_branch    <=  '1',        --  is branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write npc to register 31
                CU_writeback_mux        <=  "10"        --  write NPC
            when slli   =>
                CU_decode_ext_op        <=  "00",       --  extend as 16 bits unsigned immedaite
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "000000"    --  sll
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "01"        --  write data from ALU
            when nop    =>
                CU_decode_ext_op        <=  "00",       --  don't care
                CU_decode_dest_sel      <=  "00",       --  write to 0
                CU_decode_read1_en      <=  '0',        --  don't care
                CU_decode_read2_en      <=  '0',        --  don't care
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "000000"    --  sll
                CU_execute_top_mux      <=  '1',        --  don't care
                CU_execute_bottom_mux   <=  '1',        --  don't care
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '0',        --  don't write to rf
                CU_writeback_mux        <=  "00"        --  don't care
            when srli   =>
                CU_decode_ext_op        <=  "00",       --  extend as 16 bits unsigned immedaite
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "001000"    --  srl
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "01"        --  write data from ALU
            when srai   =>
                CU_decode_ext_op        <=  "00",       --  extend as 16 bits unsigned immedaite
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "001100"    --  sra
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "01"        --  write data from ALU
            when slti   =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immediate
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "100010"    --  slt
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "01"        --  write data from ALU
            when sgti   =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immediate
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "101010"    --  sgt
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "01"        --  write data from ALU
            when slei   =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immediate
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "100000"    --  sle
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "01"        --  write data from ALU
            when sgei   =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immediate
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "101000"    --  sge
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  don't write anything
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  '0',        --  don't care
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "01"        --  write data from ALU
            when lb     =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immediate
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "010000"    --  add
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  load
                CU_memory_signed_load   <=  '1',        --  signed load
                CU_memory_load_type     <=  "10",       --  load byte
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "00"        --  write data from MEM
            when lh     =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immediate
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "010000"    --  add
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  load
                CU_memory_signed_load   <=  '1',        --  signed load
                CU_memory_load_type     <=  "01",       --  load halfword
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "00"        --  write data from MEM
            when lw     =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immediate
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "010000"    --  add
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  load
                CU_memory_signed_load   <=  '1',        --  signed load
                CU_memory_load_type     <=  "00",       --  load word
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "00"        --  write data from MEM
            when lbu    =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immediate
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "010000"    --  add
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  load
                CU_memory_signed_load   <=  '0',        --  unsigned load
                CU_memory_load_type     <=  "10",       --  load byte
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "00"        --  write data from MEM
            when lhu    =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immediate
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "010000"    --  add
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '1',        --  load
                CU_memory_signed_load   <=  '0',        --  unsigned load
                CU_memory_load_type     <=  "01",       --  load halfword
                CU_writeback_write_en   <=  '1',        --  write to rf
                CU_writeback_mux        <=  "00"        --  write data from MEM
            when sb     =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immediate
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "010000"    --  add
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '0',        --  store
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  "01",       --  don't care
                CU_writeback_write_en   <=  '0',        --  don't write to rf
                CU_writeback_mux        <=  "00"        --  don't   --  ?
            when sh     =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immediate
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "010000"    --  add
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '0',        --  store
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  "01",       --  don't care
                CU_writeback_write_en   <=  '0',        --  don't write to rf
                CU_writeback_mux        <=  "00"        --  don't   --  ?
            when sw     =>
                CU_decode_ext_op        <=  "10",       --  extend as 16 bits signed immediate
                CU_decode_dest_sel      <=  "01",       --  use rt as destination
                CU_decode_read1_en      <=  '1',        --  read
                CU_decode_read2_en      <=  '0',        --  don't read
                CU_execute_branch_type  <=  '0',        --  don't care
                CU_execute_alu_op       <=  "010000"    --  add
                CU_execute_top_mux      <=  '1',        --  take rs
                CU_execute_bottom_mux   <=  '0',        --  read extended immediate from imm_in
                CU_execute_is_branch    <=  '0',        --  is not branch
                CU_memory_r_not_w       <=  '0',        --  store
                CU_memory_signed_load   <=  '0',        --  don't care
                CU_memory_load_type     <=  "01",       --  don't care
                CU_writeback_write_en   <=  '0',        --  don't write to rf
                CU_writeback_mux        <=  "00"        --  don't   --  ?
            when sltui  =>    --    verify if ALU supports them
            when sgtui  =>    --    verify if ALU supports them
            when sleui  =>    --    verify if ALU supports them
            when sgeui  =>    --    verify if ALU supports them
            when others =>
        end case;
    end process;

end architecture bhv;

configuration CFG_CU_CORE_BHV of cu_core is
    for bhv
    end for;
end configuration CFG_CU_CORE_BHV;
